
module reg_7 ( RST_n, VIN, d, CLK, q );
  input [13:0] d;
  output [13:0] q;
  input RST_n, VIN, CLK;
  wire   n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87;

  DFFR_X1 q_reg_4_ ( .D(n55), .CK(CLK), .RN(RST_n), .Q(q[4]), .QN(n64) );
  DFFR_X1 q_reg_3_ ( .D(n56), .CK(CLK), .RN(RST_n), .Q(q[3]), .QN(n63) );
  DFFR_X1 q_reg_2_ ( .D(n57), .CK(CLK), .RN(RST_n), .Q(q[2]), .QN(n62) );
  DFFR_X1 q_reg_1_ ( .D(n58), .CK(CLK), .RN(RST_n), .Q(q[1]), .QN(n61) );
  DFFR_X1 q_reg_0_ ( .D(n59), .CK(CLK), .RN(RST_n), .Q(q[0]), .QN(n60) );
  DFFR_X1 q_reg_5_ ( .D(n54), .CK(CLK), .RN(RST_n), .Q(q[5]), .QN(n65) );
  DFFR_X1 q_reg_6_ ( .D(n53), .CK(CLK), .RN(RST_n), .Q(q[6]), .QN(n66) );
  DFFR_X1 q_reg_7_ ( .D(n52), .CK(CLK), .RN(RST_n), .Q(q[7]), .QN(n67) );
  DFFR_X1 q_reg_8_ ( .D(n51), .CK(CLK), .RN(RST_n), .Q(q[8]), .QN(n68) );
  DFFR_X1 q_reg_9_ ( .D(n50), .CK(CLK), .RN(RST_n), .Q(q[9]), .QN(n69) );
  DFFR_X1 q_reg_10_ ( .D(n49), .CK(CLK), .RN(RST_n), .Q(q[10]), .QN(n70) );
  DFFR_X1 q_reg_11_ ( .D(n48), .CK(CLK), .RN(RST_n), .Q(q[11]), .QN(n71) );
  DFFR_X1 q_reg_12_ ( .D(n47), .CK(CLK), .RN(RST_n), .Q(q[12]), .QN(n72) );
  DFFR_X1 q_reg_13_ ( .D(n46), .CK(CLK), .RN(RST_n), .Q(q[13]), .QN(n73) );
  BUF_X1 U2 ( .A(VIN), .Z(n44) );
  BUF_X1 U3 ( .A(VIN), .Z(n43) );
  BUF_X1 U4 ( .A(VIN), .Z(n45) );
  OAI21_X1 U5 ( .B1(n44), .B2(n61), .A(n86), .ZN(n58) );
  NAND2_X1 U6 ( .A1(d[1]), .A2(n43), .ZN(n86) );
  OAI21_X1 U7 ( .B1(n44), .B2(n65), .A(n82), .ZN(n54) );
  NAND2_X1 U8 ( .A1(d[5]), .A2(n43), .ZN(n82) );
  OAI21_X1 U9 ( .B1(n44), .B2(n66), .A(n81), .ZN(n53) );
  NAND2_X1 U10 ( .A1(d[6]), .A2(n43), .ZN(n81) );
  OAI21_X1 U11 ( .B1(n44), .B2(n68), .A(n79), .ZN(n51) );
  NAND2_X1 U12 ( .A1(d[8]), .A2(n44), .ZN(n79) );
  OAI21_X1 U13 ( .B1(n44), .B2(n70), .A(n77), .ZN(n49) );
  NAND2_X1 U14 ( .A1(d[10]), .A2(n44), .ZN(n77) );
  OAI21_X1 U15 ( .B1(n44), .B2(n60), .A(n87), .ZN(n59) );
  NAND2_X1 U16 ( .A1(d[0]), .A2(n43), .ZN(n87) );
  OAI21_X1 U17 ( .B1(n44), .B2(n67), .A(n80), .ZN(n52) );
  NAND2_X1 U18 ( .A1(d[7]), .A2(n43), .ZN(n80) );
  OAI21_X1 U19 ( .B1(n44), .B2(n69), .A(n78), .ZN(n50) );
  NAND2_X1 U20 ( .A1(d[9]), .A2(n43), .ZN(n78) );
  OAI21_X1 U21 ( .B1(n44), .B2(n71), .A(n76), .ZN(n48) );
  NAND2_X1 U22 ( .A1(d[11]), .A2(n43), .ZN(n76) );
  OAI21_X1 U23 ( .B1(n44), .B2(n72), .A(n75), .ZN(n47) );
  NAND2_X1 U24 ( .A1(d[12]), .A2(n43), .ZN(n75) );
  OAI21_X1 U25 ( .B1(n44), .B2(n73), .A(n74), .ZN(n46) );
  NAND2_X1 U26 ( .A1(d[13]), .A2(n43), .ZN(n74) );
  OAI21_X1 U27 ( .B1(n45), .B2(n62), .A(n85), .ZN(n57) );
  NAND2_X1 U28 ( .A1(d[2]), .A2(n43), .ZN(n85) );
  OAI21_X1 U29 ( .B1(n45), .B2(n63), .A(n84), .ZN(n56) );
  NAND2_X1 U30 ( .A1(d[3]), .A2(n43), .ZN(n84) );
  OAI21_X1 U31 ( .B1(n45), .B2(n64), .A(n83), .ZN(n55) );
  NAND2_X1 U32 ( .A1(d[4]), .A2(n43), .ZN(n83) );
endmodule


module reg_0 ( RST_n, VIN, d, CLK, q );
  input [13:0] d;
  output [13:0] q;
  input RST_n, VIN, CLK;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  DFFR_X1 q_reg_13_ ( .D(n42), .CK(CLK), .RN(n46), .Q(q[13]), .QN(n15) );
  DFFR_X1 q_reg_12_ ( .D(n41), .CK(CLK), .RN(n46), .Q(q[12]), .QN(n16) );
  DFFR_X1 q_reg_11_ ( .D(n40), .CK(CLK), .RN(n46), .Q(q[11]), .QN(n17) );
  DFFR_X1 q_reg_10_ ( .D(n39), .CK(CLK), .RN(n46), .Q(q[10]), .QN(n18) );
  DFFR_X1 q_reg_9_ ( .D(n38), .CK(CLK), .RN(n46), .Q(q[9]), .QN(n19) );
  DFFR_X1 q_reg_8_ ( .D(n37), .CK(CLK), .RN(n46), .Q(q[8]), .QN(n20) );
  DFFR_X1 q_reg_7_ ( .D(n36), .CK(CLK), .RN(n46), .Q(q[7]), .QN(n21) );
  DFFR_X1 q_reg_6_ ( .D(n35), .CK(CLK), .RN(n46), .Q(q[6]), .QN(n22) );
  DFFR_X1 q_reg_5_ ( .D(n34), .CK(CLK), .RN(n46), .Q(q[5]), .QN(n23) );
  DFFR_X1 q_reg_4_ ( .D(n33), .CK(CLK), .RN(n46), .Q(q[4]), .QN(n24) );
  DFFR_X1 q_reg_3_ ( .D(n32), .CK(CLK), .RN(n46), .Q(q[3]), .QN(n25) );
  DFFR_X1 q_reg_2_ ( .D(n31), .CK(CLK), .RN(n46), .Q(q[2]), .QN(n26) );
  DFFR_X1 q_reg_1_ ( .D(n30), .CK(CLK), .RN(n47), .Q(q[1]), .QN(n27) );
  DFFR_X1 q_reg_0_ ( .D(n29), .CK(CLK), .RN(n47), .Q(q[0]), .QN(n28) );
  BUF_X1 U2 ( .A(VIN), .Z(n44) );
  BUF_X1 U3 ( .A(VIN), .Z(n43) );
  BUF_X1 U4 ( .A(VIN), .Z(n45) );
  BUF_X1 U5 ( .A(RST_n), .Z(n46) );
  BUF_X1 U6 ( .A(RST_n), .Z(n47) );
  OAI21_X1 U7 ( .B1(n44), .B2(n28), .A(n1), .ZN(n29) );
  NAND2_X1 U8 ( .A1(d[0]), .A2(n43), .ZN(n1) );
  OAI21_X1 U9 ( .B1(n44), .B2(n27), .A(n2), .ZN(n30) );
  NAND2_X1 U10 ( .A1(d[1]), .A2(n43), .ZN(n2) );
  OAI21_X1 U11 ( .B1(n44), .B2(n23), .A(n6), .ZN(n34) );
  NAND2_X1 U12 ( .A1(d[5]), .A2(n43), .ZN(n6) );
  OAI21_X1 U13 ( .B1(n44), .B2(n22), .A(n7), .ZN(n35) );
  NAND2_X1 U14 ( .A1(d[6]), .A2(n43), .ZN(n7) );
  OAI21_X1 U15 ( .B1(n44), .B2(n21), .A(n8), .ZN(n36) );
  NAND2_X1 U16 ( .A1(d[7]), .A2(n43), .ZN(n8) );
  OAI21_X1 U17 ( .B1(n44), .B2(n19), .A(n10), .ZN(n38) );
  NAND2_X1 U18 ( .A1(d[9]), .A2(n43), .ZN(n10) );
  OAI21_X1 U19 ( .B1(n44), .B2(n17), .A(n12), .ZN(n40) );
  NAND2_X1 U20 ( .A1(d[11]), .A2(n43), .ZN(n12) );
  OAI21_X1 U21 ( .B1(n44), .B2(n16), .A(n13), .ZN(n41) );
  NAND2_X1 U22 ( .A1(d[12]), .A2(n43), .ZN(n13) );
  OAI21_X1 U23 ( .B1(n44), .B2(n15), .A(n14), .ZN(n42) );
  NAND2_X1 U24 ( .A1(d[13]), .A2(n43), .ZN(n14) );
  OAI21_X1 U25 ( .B1(n44), .B2(n20), .A(n9), .ZN(n37) );
  NAND2_X1 U26 ( .A1(d[8]), .A2(n44), .ZN(n9) );
  OAI21_X1 U27 ( .B1(n44), .B2(n18), .A(n11), .ZN(n39) );
  NAND2_X1 U28 ( .A1(d[10]), .A2(n44), .ZN(n11) );
  OAI21_X1 U29 ( .B1(n45), .B2(n26), .A(n3), .ZN(n31) );
  NAND2_X1 U30 ( .A1(d[2]), .A2(n43), .ZN(n3) );
  OAI21_X1 U31 ( .B1(n45), .B2(n25), .A(n4), .ZN(n32) );
  NAND2_X1 U32 ( .A1(d[3]), .A2(n43), .ZN(n4) );
  OAI21_X1 U33 ( .B1(n45), .B2(n24), .A(n5), .ZN(n33) );
  NAND2_X1 U34 ( .A1(d[4]), .A2(n43), .ZN(n5) );
endmodule


module IIR_ADV ( CLK, RST_n, VIN, DIN, B0, B1, B2, B3, A1, A2, VOUT, DOUT );
  input [13:0] DIN;
  input [13:0] B0;
  input [13:0] B1;
  input [13:0] B2;
  input [13:0] B3;
  input [13:0] A1;
  input [13:0] A2;
  output [13:0] DOUT;
  input CLK, RST_n, VIN;
  output VOUT;
  wire   n185, n30, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, REGISTER1_n266, REGISTER1_n265, REGISTER1_n264,
         REGISTER1_n263, REGISTER1_n262, REGISTER1_n261, REGISTER1_n260,
         REGISTER1_n259, REGISTER1_n258, REGISTER1_n257, REGISTER1_n256,
         REGISTER1_n255, REGISTER1_n254, REGISTER1_n253, REG1_1_n267,
         REG1_1_n266, REG1_1_n265, REG1_1_n264, REG1_1_n263, REG1_1_n262,
         REG1_1_n261, REG1_1_n260, REG1_1_n259, REG1_1_n258, REG1_1_n257,
         REG1_1_n256, REG1_1_n255, REG1_1_n254, REGISTER2_n266, REGISTER2_n265,
         REGISTER2_n264, REGISTER2_n263, REGISTER2_n262, REGISTER2_n261,
         REGISTER2_n260, REGISTER2_n259, REGISTER2_n258, REGISTER2_n257,
         REGISTER2_n256, REGISTER2_n255, REGISTER2_n254, REGISTER2_n253,
         REG2_1_n272, REG2_1_n271, REG2_1_n92, REG2_1_n75, REG2_1_n270,
         REG2_1_n269, REG2_1_n268, REG2_1_n267, REG2_1_n266, REG2_1_n265,
         REG2_1_n264, REG2_1_n263, REG2_1_n262, REG2_1_n261, REG2_1_n260,
         REG2_1_n259, REG2_1_n258, REGISTER3_n266, REGISTER3_n265,
         REGISTER3_n264, REGISTER3_n263, REGISTER3_n262, REGISTER3_n261,
         REGISTER3_n260, REGISTER3_n259, REGISTER3_n258, REGISTER3_n257,
         REGISTER3_n256, REGISTER3_n255, REGISTER3_n254, REGISTER3_n253,
         REG3_1_n267, REG3_1_n266, REG3_1_n265, REG3_1_n264, REG3_1_n263,
         REG3_1_n262, REG3_1_n261, REG3_1_n260, REG3_1_n259, REG3_1_n258,
         REG3_1_n257, REG3_1_n256, REG3_1_n255, REG3_1_n254, REGISTER4_n266,
         REGISTER4_n265, REGISTER4_n264, REGISTER4_n263, REGISTER4_n262,
         REGISTER4_n261, REGISTER4_n260, REGISTER4_n259, REGISTER4_n258,
         REGISTER4_n257, REGISTER4_n256, REGISTER4_n255, REGISTER4_n254,
         REGISTER4_n253, REG4_1_n266, REG4_1_n265, REG4_1_n264, REG4_1_n263,
         REG4_1_n262, REG4_1_n261, REG4_1_n260, REG4_1_n259, REG4_1_n258,
         REG4_1_n257, REG4_1_n256, REG4_1_n255, REG4_1_n254, REG4_1_n253,
         SUB1_N1, SUB1_N10, SUB1_N11, SUB1_N12, SUB1_N13, SUB1_N2, SUB1_N3,
         SUB1_N4, SUB1_N5, SUB1_N6, SUB1_N7, SUB1_N8, SUB1_N9, REG11_n64,
         REG11_n266, REG11_n265, REG11_n264, REG11_n263, REG11_n262,
         REG11_n261, REG11_n260, REG11_n259, REG11_n258, REG11_n257,
         REG11_n256, REG11_n255, REG11_n254, REG21_n266, REG21_n265,
         REG21_n264, REG21_n263, REG21_n262, REG21_n261, REG21_n260,
         REG21_n259, REG21_n258, REG21_n257, REG21_n256, REG21_n255,
         REG21_n254, REG21_n253, REG31_n266, REG31_n265, REG31_n264,
         REG31_n263, REG31_n262, REG31_n261, REG31_n260, REG31_n259,
         REG31_n258, REG31_n257, REG31_n256, REG31_n255, REG31_n254,
         REG31_n253, REG41_n266, REG41_n265, REG41_n264, REG41_n263,
         REG41_n262, REG41_n261, REG41_n260, REG41_n259, REG41_n258,
         REG41_n257, REG41_n256, REG41_n255, REG41_n254, REG41_n253,
         REG51_n266, REG51_n265, REG51_n264, REG51_n263, REG51_n262,
         REG51_n261, REG51_n260, REG51_n259, REG51_n258, REG51_n257,
         REG51_n256, REG51_n255, REG51_n254, REG51_n253, REG61_n267,
         REG61_n266, REG61_n265, REG61_n264, REG61_n263, REG61_n262,
         REG61_n261, REG61_n260, REG61_n259, REG61_n258, REG61_n257,
         REG61_n256, REG61_n255, REG61_n254, sig_ff2_9_, sig_ff2_8_,
         sig_ff2_7_, sig_ff2_6_, sig_ff2_5_, sig_ff2_4_, sig_ff2_3_,
         sig_ff2_2_, sig_ff2_1_, sig_ff2_13_, sig_ff2_12_, sig_ff2_11_,
         sig_ff2_10_, sig_ff2_0_, sig_ff1_9_, sig_ff1_8_, sig_ff1_7_,
         sig_ff1_6_, sig_ff1_5_, sig_ff1_4_, sig_ff1_3_, sig_ff1_2_,
         sig_ff1_1_, sig_ff1_13_, sig_ff1_12_, sig_ff1_11_, sig_ff1_10_,
         sig_ff1_0_, fb_9_, fb_8_, fb_7_, fb_6_, fb_5_, fb_4_, fb_3_, fb_2_,
         fb_1_, fb_13_, fb_12_, fb_11_, fb_10_, fb_0_, n259, n260, n262, n263,
         n264, n266, n267, n268, n269, n271, n272, n273, n274, n276, n277,
         n278, n279, n280, n282, n283, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, p6_mult_21_n844, p6_mult_21_n843, p6_mult_21_n842,
         p6_mult_21_n841, p6_mult_21_n840, p6_mult_21_n839, p6_mult_21_n838,
         p6_mult_21_n837, p6_mult_21_n831, p6_mult_21_n830, p6_mult_21_n829,
         p6_mult_21_n828, p6_mult_21_n827, p6_mult_21_n826, p6_mult_21_n825,
         p6_mult_21_n824, p6_mult_21_n823, p6_mult_21_n822, p6_mult_21_n821,
         p6_mult_21_n820, p6_mult_21_n819, p6_mult_21_n818, p6_mult_21_n817,
         p6_mult_21_n816, p6_mult_21_n815, p6_mult_21_n813, p6_mult_21_n811,
         p6_mult_21_n809, p6_mult_21_n808, p6_mult_21_n807, p6_mult_21_n806,
         p6_mult_21_n805, p6_mult_21_n804, p6_mult_21_n803, p6_mult_21_n802,
         p6_mult_21_n801, p6_mult_21_n800, p6_mult_21_n799, p6_mult_21_n798,
         p6_mult_21_n797, p6_mult_21_n796, p6_mult_21_n795, p6_mult_21_n794,
         p6_mult_21_n793, p6_mult_21_n792, p6_mult_21_n791, p6_mult_21_n790,
         p6_mult_21_n789, p6_mult_21_n788, p6_mult_21_n787, p6_mult_21_n786,
         p6_mult_21_n785, p6_mult_21_n784, p6_mult_21_n783, p6_mult_21_n782,
         p6_mult_21_n781, p6_mult_21_n780, p6_mult_21_n779, p6_mult_21_n778,
         p6_mult_21_n777, p6_mult_21_n776, p6_mult_21_n774, p6_mult_21_n773,
         p6_mult_21_n772, p6_mult_21_n771, p6_mult_21_n770, p6_mult_21_n769,
         p6_mult_21_n768, p6_mult_21_n767, p6_mult_21_n766, p6_mult_21_n765,
         p6_mult_21_n764, p6_mult_21_n763, p6_mult_21_n762, p6_mult_21_n761,
         p6_mult_21_n760, p6_mult_21_n759, p6_mult_21_n757, p6_mult_21_n756,
         p6_mult_21_n755, p6_mult_21_n754, p6_mult_21_n753, p6_mult_21_n752,
         p6_mult_21_n751, p6_mult_21_n750, p6_mult_21_n749, p6_mult_21_n748,
         p6_mult_21_n747, p6_mult_21_n746, p6_mult_21_n745, p6_mult_21_n744,
         p6_mult_21_n743, p6_mult_21_n742, p6_mult_21_n740, p6_mult_21_n739,
         p6_mult_21_n738, p6_mult_21_n737, p6_mult_21_n736, p6_mult_21_n735,
         p6_mult_21_n734, p6_mult_21_n733, p6_mult_21_n732, p6_mult_21_n731,
         p6_mult_21_n730, p6_mult_21_n729, p6_mult_21_n728, p6_mult_21_n727,
         p6_mult_21_n726, p6_mult_21_n725, p6_mult_21_n724, p6_mult_21_n723,
         p6_mult_21_n722, p6_mult_21_n721, p6_mult_21_n720, p6_mult_21_n719,
         p6_mult_21_n718, p6_mult_21_n717, p6_mult_21_n716, p6_mult_21_n715,
         p6_mult_21_n714, p6_mult_21_n713, p6_mult_21_n712, p6_mult_21_n711,
         p6_mult_21_n710, p6_mult_21_n709, p6_mult_21_n708, p6_mult_21_n707,
         p6_mult_21_n706, p6_mult_21_n705, p6_mult_21_n704, p6_mult_21_n703,
         p6_mult_21_n702, p6_mult_21_n701, p6_mult_21_n700, p6_mult_21_n699,
         p6_mult_21_n698, p6_mult_21_n697, p6_mult_21_n696, p6_mult_21_n695,
         p6_mult_21_n694, p6_mult_21_n693, p6_mult_21_n692, p6_mult_21_n691,
         p6_mult_21_n690, p6_mult_21_n689, p6_mult_21_n688, p6_mult_21_n687,
         p6_mult_21_n686, p6_mult_21_n681, p6_mult_21_n680, p6_mult_21_n679,
         p6_mult_21_n678, p6_mult_21_n674, p6_mult_21_n673, p6_mult_21_n672,
         p6_mult_21_n671, p6_mult_21_n667, p6_mult_21_n661, p6_mult_21_n660,
         p6_mult_21_n659, p6_mult_21_n651, p6_mult_21_n647, p6_mult_21_n643,
         p6_mult_21_n642, p6_mult_21_n641, p6_mult_21_n640, p6_mult_21_n636,
         p6_mult_21_n635, p6_mult_21_n418, p6_mult_21_n417, p6_mult_21_n416,
         p6_mult_21_n415, p6_mult_21_n414, p6_mult_21_n413, p6_mult_21_n412,
         p6_mult_21_n411, p6_mult_21_n410, p6_mult_21_n409, p6_mult_21_n408,
         p6_mult_21_n405, p6_mult_21_n404, p6_mult_21_n403, p6_mult_21_n402,
         p6_mult_21_n401, p6_mult_21_n400, p6_mult_21_n399, p6_mult_21_n398,
         p6_mult_21_n397, p6_mult_21_n396, p6_mult_21_n395, p6_mult_21_n394,
         p6_mult_21_n393, p6_mult_21_n392, p6_mult_21_n390, p6_mult_21_n389,
         p6_mult_21_n388, p6_mult_21_n387, p6_mult_21_n386, p6_mult_21_n385,
         p6_mult_21_n384, p6_mult_21_n382, p6_mult_21_n381, p6_mult_21_n380,
         p6_mult_21_n379, p6_mult_21_n377, p6_mult_21_n376, p6_mult_21_n375,
         p6_mult_21_n374, p6_mult_21_n373, p6_mult_21_n372, p6_mult_21_n371,
         p6_mult_21_n370, p6_mult_21_n369, p6_mult_21_n368, p6_mult_21_n367,
         p6_mult_21_n366, p6_mult_21_n365, p6_mult_21_n363, p6_mult_21_n362,
         p6_mult_21_n361, p6_mult_21_n360, p6_mult_21_n359, p6_mult_21_n358,
         p6_mult_21_n357, p6_mult_21_n356, p6_mult_21_n355, p6_mult_21_n354,
         p6_mult_21_n353, p6_mult_21_n352, p6_mult_21_n351, p6_mult_21_n349,
         p6_mult_21_n348, p6_mult_21_n346, p6_mult_21_n345, p6_mult_21_n344,
         p6_mult_21_n343, p6_mult_21_n342, p6_mult_21_n341, p6_mult_21_n340,
         p6_mult_21_n339, p6_mult_21_n338, p6_mult_21_n337, p6_mult_21_n336,
         p6_mult_21_n335, p6_mult_21_n334, p6_mult_21_n333, p6_mult_21_n332,
         p6_mult_21_n331, p6_mult_21_n330, p6_mult_21_n329, p6_mult_21_n328,
         p6_mult_21_n327, p6_mult_21_n326, p6_mult_21_n325, p6_mult_21_n321,
         p6_mult_21_n317, p6_mult_21_n314, p6_mult_21_n313, p6_mult_21_n312,
         p6_mult_21_n311, p6_mult_21_n308, p6_mult_21_n307, p6_mult_21_n304,
         p6_mult_21_n303, p6_mult_21_n302, p6_mult_21_n301, p6_mult_21_n300,
         p6_mult_21_n299, p6_mult_21_n298, p6_mult_21_n297, p6_mult_21_n296,
         p6_mult_21_n295, p6_mult_21_n294, p6_mult_21_n293, p6_mult_21_n292,
         p6_mult_21_n291, p6_mult_21_n290, p6_mult_21_n289, p6_mult_21_n288,
         p6_mult_21_n287, p6_mult_21_n286, p6_mult_21_n285, p6_mult_21_n284,
         p6_mult_21_n283, p6_mult_21_n282, p6_mult_21_n281, p6_mult_21_n280,
         p6_mult_21_n279, p6_mult_21_n278, p6_mult_21_n277, p6_mult_21_n276,
         p6_mult_21_n275, p6_mult_21_n274, p6_mult_21_n273, p6_mult_21_n272,
         p6_mult_21_n271, p6_mult_21_n270, p6_mult_21_n269, p6_mult_21_n268,
         p6_mult_21_n267, p6_mult_21_n266, p6_mult_21_n265, p6_mult_21_n264,
         p6_mult_21_n263, p6_mult_21_n262, p6_mult_21_n261, p6_mult_21_n260,
         p6_mult_21_n259, p6_mult_21_n258, p6_mult_21_n257, p6_mult_21_n256,
         p6_mult_21_n255, p6_mult_21_n254, p6_mult_21_n253, p6_mult_21_n252,
         p6_mult_21_n251, p6_mult_21_n250, p6_mult_21_n249, p6_mult_21_n248,
         p6_mult_21_n247, p6_mult_21_n246, p6_mult_21_n245, p6_mult_21_n244,
         p6_mult_21_n243, p6_mult_21_n242, p6_mult_21_n241, p6_mult_21_n240,
         p6_mult_21_n239, p6_mult_21_n238, p6_mult_21_n237, p6_mult_21_n236,
         p6_mult_21_n235, p6_mult_21_n234, p6_mult_21_n233, p6_mult_21_n232,
         p6_mult_21_n231, p6_mult_21_n230, p6_mult_21_n229, p6_mult_21_n228,
         p6_mult_21_n227, p6_mult_21_n226, p6_mult_21_n225, p6_mult_21_n224,
         p6_mult_21_n223, p6_mult_21_n222, p6_mult_21_n221, p6_mult_21_n220,
         p6_mult_21_n219, p6_mult_21_n218, p6_mult_21_n217, p6_mult_21_n216,
         p6_mult_21_n215, p6_mult_21_n214, p6_mult_21_n213, p6_mult_21_n212,
         p6_mult_21_n211, p6_mult_21_n210, p6_mult_21_n209, p6_mult_21_n208,
         p6_mult_21_n207, p6_mult_21_n206, p6_mult_21_n205, p6_mult_21_n204,
         p6_mult_21_n203, p6_mult_21_n202, p6_mult_21_n201, p6_mult_21_n200,
         p6_mult_21_n199, p6_mult_21_n198, p6_mult_21_n197, p6_mult_21_n196,
         p6_mult_21_n195, p6_mult_21_n194, p6_mult_21_n193, p6_mult_21_n192,
         p6_mult_21_n191, p6_mult_21_n190, p6_mult_21_n189, p6_mult_21_n188,
         p6_mult_21_n187, p6_mult_21_n186, p6_mult_21_n185, p6_mult_21_n184,
         p6_mult_21_n183, p6_mult_21_n182, p6_mult_21_n181, p6_mult_21_n180,
         p6_mult_21_n179, p6_mult_21_n178, p6_mult_21_n177, p6_mult_21_n176,
         p6_mult_21_n175, p6_mult_21_n174, p6_mult_21_n173, p6_mult_21_n172,
         p6_mult_21_n171, p6_mult_21_n170, p6_mult_21_n169, p6_mult_21_n168,
         p6_mult_21_n167, p6_mult_21_n166, p6_mult_21_n165, p6_mult_21_n164,
         p6_mult_21_n163, p6_mult_21_n162, p6_mult_21_n149, p6_mult_21_n148,
         p6_mult_21_n147, p6_mult_21_n146, p6_mult_21_n145, p6_mult_21_n144,
         p6_mult_21_n143, p6_mult_21_n142, p6_mult_21_n141, p6_mult_21_n140,
         p6_mult_21_n139, p6_mult_21_n138, p6_mult_21_n137, p6_mult_21_n136,
         p7_mult_21_n1034, p7_mult_21_n1404, p7_mult_21_n1403,
         p7_mult_21_n1402, p7_mult_21_n1401, p7_mult_21_n1400,
         p7_mult_21_n1399, p7_mult_21_n1398, p7_mult_21_n1397,
         p7_mult_21_n1396, p7_mult_21_n1395, p7_mult_21_n1394,
         p7_mult_21_n1393, p7_mult_21_n1392, p7_mult_21_n1391,
         p7_mult_21_n1390, p7_mult_21_n1389, p7_mult_21_n1388,
         p7_mult_21_n1387, p7_mult_21_n1386, p7_mult_21_n1385,
         p7_mult_21_n1384, p7_mult_21_n1383, p7_mult_21_n1382,
         p7_mult_21_n1381, p7_mult_21_n1380, p7_mult_21_n1379,
         p7_mult_21_n1378, p7_mult_21_n1377, p7_mult_21_n1376,
         p7_mult_21_n1375, p7_mult_21_n1374, p7_mult_21_n1373,
         p7_mult_21_n1372, p7_mult_21_n1371, p7_mult_21_n1370,
         p7_mult_21_n1369, p7_mult_21_n1368, p7_mult_21_n1367,
         p7_mult_21_n1366, p7_mult_21_n1365, p7_mult_21_n1364,
         p7_mult_21_n1363, p7_mult_21_n1362, p7_mult_21_n1361,
         p7_mult_21_n1360, p7_mult_21_n1359, p7_mult_21_n1358,
         p7_mult_21_n1357, p7_mult_21_n1356, p7_mult_21_n1355,
         p7_mult_21_n1354, p7_mult_21_n1353, p7_mult_21_n1352,
         p7_mult_21_n1351, p7_mult_21_n1350, p7_mult_21_n1348,
         p7_mult_21_n1347, p7_mult_21_n1346, p7_mult_21_n1345,
         p7_mult_21_n1344, p7_mult_21_n1343, p7_mult_21_n1342,
         p7_mult_21_n1341, p7_mult_21_n1340, p7_mult_21_n1339,
         p7_mult_21_n1338, p7_mult_21_n1337, p7_mult_21_n1336,
         p7_mult_21_n1335, p7_mult_21_n1333, p7_mult_21_n1332,
         p7_mult_21_n1331, p7_mult_21_n1329, p7_mult_21_n1328,
         p7_mult_21_n1327, p7_mult_21_n1326, p7_mult_21_n1325,
         p7_mult_21_n1324, p7_mult_21_n1323, p7_mult_21_n1322,
         p7_mult_21_n1321, p7_mult_21_n1320, p7_mult_21_n1319,
         p7_mult_21_n1318, p7_mult_21_n1317, p7_mult_21_n1316,
         p7_mult_21_n1315, p7_mult_21_n1314, p7_mult_21_n1313,
         p7_mult_21_n1312, p7_mult_21_n1311, p7_mult_21_n1310,
         p7_mult_21_n1308, p7_mult_21_n1307, p7_mult_21_n1305,
         p7_mult_21_n1304, p7_mult_21_n1303, p7_mult_21_n1302,
         p7_mult_21_n1301, p7_mult_21_n1300, p7_mult_21_n1299,
         p7_mult_21_n1298, p7_mult_21_n1297, p7_mult_21_n1296,
         p7_mult_21_n1295, p7_mult_21_n1294, p7_mult_21_n1293,
         p7_mult_21_n1292, p7_mult_21_n1291, p7_mult_21_n1290,
         p7_mult_21_n1289, p7_mult_21_n1288, p7_mult_21_n1287,
         p7_mult_21_n1286, p7_mult_21_n1285, p7_mult_21_n1284,
         p7_mult_21_n1283, p7_mult_21_n1281, p7_mult_21_n1280,
         p7_mult_21_n1279, p7_mult_21_n1278, p7_mult_21_n1277,
         p7_mult_21_n1274, p7_mult_21_n1273, p7_mult_21_n1272,
         p7_mult_21_n1271, p7_mult_21_n1270, p7_mult_21_n1269,
         p7_mult_21_n1268, p7_mult_21_n1267, p7_mult_21_n1266,
         p7_mult_21_n1265, p7_mult_21_n1264, p7_mult_21_n1262,
         p7_mult_21_n1261, p7_mult_21_n1260, p7_mult_21_n1258,
         p7_mult_21_n1257, p7_mult_21_n1256, p7_mult_21_n1255,
         p7_mult_21_n1254, p7_mult_21_n1253, p7_mult_21_n1252,
         p7_mult_21_n1251, p7_mult_21_n1250, p7_mult_21_n1248,
         p7_mult_21_n1247, p7_mult_21_n1246, p7_mult_21_n1245,
         p7_mult_21_n1244, p7_mult_21_n1243, p7_mult_21_n1242,
         p7_mult_21_n1241, p7_mult_21_n1240, p7_mult_21_n1239,
         p7_mult_21_n1238, p7_mult_21_n1237, p7_mult_21_n1236,
         p7_mult_21_n1235, p7_mult_21_n1234, p7_mult_21_n1233,
         p7_mult_21_n1232, p7_mult_21_n1231, p7_mult_21_n1230,
         p7_mult_21_n1229, p7_mult_21_n1228, p7_mult_21_n1227,
         p7_mult_21_n1226, p7_mult_21_n1225, p7_mult_21_n1224,
         p7_mult_21_n1223, p7_mult_21_n1222, p7_mult_21_n1221,
         p7_mult_21_n1220, p7_mult_21_n1219, p7_mult_21_n1218,
         p7_mult_21_n1217, p7_mult_21_n1216, p7_mult_21_n1215,
         p7_mult_21_n1214, p7_mult_21_n1213, p7_mult_21_n1212,
         p7_mult_21_n1211, p7_mult_21_n1210, p7_mult_21_n1209,
         p7_mult_21_n1208, p7_mult_21_n1207, p7_mult_21_n1206,
         p7_mult_21_n1205, p7_mult_21_n1204, p7_mult_21_n1203,
         p7_mult_21_n1202, p7_mult_21_n1201, p7_mult_21_n1200,
         p7_mult_21_n1199, p7_mult_21_n1198, p7_mult_21_n1197,
         p7_mult_21_n1196, p7_mult_21_n1195, p7_mult_21_n1194,
         p7_mult_21_n1193, p7_mult_21_n1192, p7_mult_21_n1191,
         p7_mult_21_n1190, p7_mult_21_n1189, p7_mult_21_n1188,
         p7_mult_21_n1187, p7_mult_21_n1186, p7_mult_21_n1185,
         p7_mult_21_n1184, p7_mult_21_n1183, p7_mult_21_n1182,
         p7_mult_21_n1181, p7_mult_21_n1180, p7_mult_21_n1179,
         p7_mult_21_n1178, p7_mult_21_n1177, p7_mult_21_n1176,
         p7_mult_21_n1175, p7_mult_21_n1174, p7_mult_21_n1173,
         p7_mult_21_n1172, p7_mult_21_n1171, p7_mult_21_n1170,
         p7_mult_21_n1169, p7_mult_21_n1168, p7_mult_21_n1167,
         p7_mult_21_n1166, p7_mult_21_n1165, p7_mult_21_n1164,
         p7_mult_21_n1163, p7_mult_21_n1162, p7_mult_21_n1161,
         p7_mult_21_n1160, p7_mult_21_n1159, p7_mult_21_n1158,
         p7_mult_21_n1157, p7_mult_21_n1156, p7_mult_21_n1155,
         p7_mult_21_n1154, p7_mult_21_n1153, p7_mult_21_n1152,
         p7_mult_21_n1151, p7_mult_21_n1150, p7_mult_21_n1149,
         p7_mult_21_n1148, p7_mult_21_n1147, p7_mult_21_n1146,
         p7_mult_21_n1145, p7_mult_21_n1144, p7_mult_21_n1143,
         p7_mult_21_n1142, p7_mult_21_n1141, p7_mult_21_n1140,
         p7_mult_21_n1139, p7_mult_21_n1138, p7_mult_21_n1137,
         p7_mult_21_n1136, p7_mult_21_n1135, p7_mult_21_n1134,
         p7_mult_21_n1133, p7_mult_21_n1132, p7_mult_21_n1131,
         p7_mult_21_n1130, p7_mult_21_n1129, p7_mult_21_n1128,
         p7_mult_21_n1127, p7_mult_21_n1126, p7_mult_21_n1125,
         p7_mult_21_n1124, p7_mult_21_n1123, p7_mult_21_n1122,
         p7_mult_21_n1121, p7_mult_21_n1120, p7_mult_21_n1119,
         p7_mult_21_n1118, p7_mult_21_n1117, p7_mult_21_n1116,
         p7_mult_21_n1115, p7_mult_21_n1114, p7_mult_21_n1113,
         p7_mult_21_n1112, p7_mult_21_n1111, p7_mult_21_n1110,
         p7_mult_21_n1108, p7_mult_21_n1107, p7_mult_21_n1106,
         p7_mult_21_n1105, p7_mult_21_n1104, p7_mult_21_n1103,
         p7_mult_21_n1102, p7_mult_21_n1101, p7_mult_21_n1099,
         p7_mult_21_n1098, p7_mult_21_n1097, p7_mult_21_n1096,
         p7_mult_21_n1095, p7_mult_21_n1094, p7_mult_21_n1093,
         p7_mult_21_n1092, p7_mult_21_n1091, p7_mult_21_n1090,
         p7_mult_21_n1089, p7_mult_21_n1088, p7_mult_21_n1087,
         p7_mult_21_n1086, p7_mult_21_n1085, p7_mult_21_n1084,
         p7_mult_21_n1083, p7_mult_21_n1082, p7_mult_21_n1081,
         p7_mult_21_n1080, p7_mult_21_n1079, p7_mult_21_n1078,
         p7_mult_21_n1077, p7_mult_21_n1076, p7_mult_21_n1075,
         p7_mult_21_n1074, p7_mult_21_n1073, p7_mult_21_n1072,
         p7_mult_21_n1071, p7_mult_21_n1070, p7_mult_21_n1069,
         p7_mult_21_n1068, p7_mult_21_n1067, p7_mult_21_n1066,
         p7_mult_21_n1065, p7_mult_21_n1064, p7_mult_21_n1063,
         p7_mult_21_n1062, p7_mult_21_n1061, p7_mult_21_n1060,
         p7_mult_21_n1059, p7_mult_21_n1058, p7_mult_21_n1057,
         p7_mult_21_n1056, p7_mult_21_n1055, p7_mult_21_n1054,
         p7_mult_21_n1053, p7_mult_21_n1052, p7_mult_21_n1051,
         p7_mult_21_n1050, p7_mult_21_n1049, p7_mult_21_n1048,
         p7_mult_21_n1047, p7_mult_21_n1046, p7_mult_21_n1045,
         p7_mult_21_n1044, p7_mult_21_n1043, p7_mult_21_n1042,
         p7_mult_21_n1041, p7_mult_21_n1040, p7_mult_21_n1039,
         p7_mult_21_n1038, p7_mult_21_n1037, p7_mult_21_n1036,
         p7_mult_21_n1035, p7_mult_21_n1033, p7_mult_21_n1032,
         p7_mult_21_n1031, p7_mult_21_n1030, p7_mult_21_n1029,
         p7_mult_21_n1028, p7_mult_21_n1027, p7_mult_21_n1026,
         p7_mult_21_n1025, p7_mult_21_n1024, p7_mult_21_n1023,
         p7_mult_21_n1022, p7_mult_21_n1021, p7_mult_21_n1020,
         p7_mult_21_n1019, p7_mult_21_n1018, p7_mult_21_n1017,
         p7_mult_21_n1016, p7_mult_21_n1015, p7_mult_21_n1014,
         p7_mult_21_n1013, p7_mult_21_n1012, p7_mult_21_n1011,
         p7_mult_21_n1010, p7_mult_21_n1009, p7_mult_21_n1008,
         p7_mult_21_n1007, p7_mult_21_n1006, p7_mult_21_n1005,
         p7_mult_21_n1004, p7_mult_21_n1003, p7_mult_21_n1002,
         p7_mult_21_n1001, p7_mult_21_n1000, p7_mult_21_n999, p7_mult_21_n998,
         p7_mult_21_n997, p7_mult_21_n996, p7_mult_21_n995, p7_mult_21_n994,
         p7_mult_21_n993, p7_mult_21_n992, p7_mult_21_n991, p7_mult_21_n990,
         p7_mult_21_n989, p7_mult_21_n988, p7_mult_21_n987, p7_mult_21_n986,
         p7_mult_21_n985, p7_mult_21_n984, p7_mult_21_n983, p7_mult_21_n982,
         p7_mult_21_n981, p7_mult_21_n980, p7_mult_21_n979, p7_mult_21_n978,
         p7_mult_21_n977, p7_mult_21_n976, p7_mult_21_n975, p7_mult_21_n974,
         p7_mult_21_n972, p7_mult_21_n971, p7_mult_21_n970, p7_mult_21_n969,
         p7_mult_21_n968, p7_mult_21_n967, p7_mult_21_n966, p7_mult_21_n965,
         p7_mult_21_n964, p7_mult_21_n963, p7_mult_21_n962, p7_mult_21_n961,
         p7_mult_21_n960, p7_mult_21_n959, p7_mult_21_n958, p7_mult_21_n957,
         p7_mult_21_n956, p7_mult_21_n955, p7_mult_21_n954, p7_mult_21_n953,
         p7_mult_21_n952, p7_mult_21_n951, p7_mult_21_n950, p7_mult_21_n949,
         p7_mult_21_n948, p7_mult_21_n947, p7_mult_21_n946, p7_mult_21_n945,
         p7_mult_21_n944, p7_mult_21_n943, p7_mult_21_n942, p7_mult_21_n941,
         p7_mult_21_n940, p7_mult_21_n939, p7_mult_21_n938, p7_mult_21_n937,
         p7_mult_21_n936, p7_mult_21_n935, p7_mult_21_n934, p7_mult_21_n933,
         p7_mult_21_n932, p7_mult_21_n931, p7_mult_21_n930, p7_mult_21_n929,
         p7_mult_21_n928, p7_mult_21_n927, p7_mult_21_n926, p7_mult_21_n925,
         p7_mult_21_n924, p7_mult_21_n923, p7_mult_21_n922, p7_mult_21_n921,
         p7_mult_21_n920, p7_mult_21_n919, p7_mult_21_n918, p7_mult_21_n917,
         p7_mult_21_n916, p7_mult_21_n915, p7_mult_21_n914, p7_mult_21_n913,
         p7_mult_21_n912, p7_mult_21_n911, p7_mult_21_n910, p7_mult_21_n909,
         p7_mult_21_n908, p7_mult_21_n907, p7_mult_21_n906, p7_mult_21_n905,
         p7_mult_21_n904, p7_mult_21_n903, p7_mult_21_n902, p7_mult_21_n901,
         p7_mult_21_n900, p7_mult_21_n899, p7_mult_21_n898, p7_mult_21_n897,
         p7_mult_21_n896, p7_mult_21_n895, p7_mult_21_n894, p7_mult_21_n893,
         p7_mult_21_n892, p7_mult_21_n891, p7_mult_21_n890, p7_mult_21_n889,
         p7_mult_21_n888, p7_mult_21_n887, p7_mult_21_n886, p7_mult_21_n885,
         p7_mult_21_n884, p7_mult_21_n883, p7_mult_21_n882, p7_mult_21_n880,
         p7_mult_21_n878, p7_mult_21_n877, p7_mult_21_n876, p7_mult_21_n875,
         p7_mult_21_n874, p7_mult_21_n873, p7_mult_21_n872, p7_mult_21_n871,
         p7_mult_21_n870, p7_mult_21_n869, p7_mult_21_n868, p7_mult_21_n867,
         p7_mult_21_n866, p7_mult_21_n865, p7_mult_21_n864, p7_mult_21_n860,
         p7_mult_21_n852, p7_mult_21_n847, p7_mult_21_n846, p7_mult_21_n844,
         p8_mult_21_n837, p8_mult_21_n836, p8_mult_21_n832, p8_mult_21_n826,
         p8_mult_21_n825, p8_mult_21_n824, p8_mult_21_n823, p8_mult_21_n822,
         p8_mult_21_n821, p8_mult_21_n820, p8_mult_21_n819, p8_mult_21_n818,
         p8_mult_21_n817, p8_mult_21_n816, p8_mult_21_n815, p8_mult_21_n814,
         p8_mult_21_n812, p8_mult_21_n810, p8_mult_21_n808, p8_mult_21_n806,
         p8_mult_21_n805, p8_mult_21_n804, p8_mult_21_n803, p8_mult_21_n802,
         p8_mult_21_n801, p8_mult_21_n800, p8_mult_21_n799, p8_mult_21_n798,
         p8_mult_21_n797, p8_mult_21_n796, p8_mult_21_n795, p8_mult_21_n794,
         p8_mult_21_n793, p8_mult_21_n792, p8_mult_21_n791, p8_mult_21_n790,
         p8_mult_21_n789, p8_mult_21_n788, p8_mult_21_n787, p8_mult_21_n786,
         p8_mult_21_n785, p8_mult_21_n784, p8_mult_21_n783, p8_mult_21_n782,
         p8_mult_21_n781, p8_mult_21_n780, p8_mult_21_n779, p8_mult_21_n778,
         p8_mult_21_n777, p8_mult_21_n776, p8_mult_21_n775, p8_mult_21_n773,
         p8_mult_21_n772, p8_mult_21_n771, p8_mult_21_n770, p8_mult_21_n769,
         p8_mult_21_n768, p8_mult_21_n767, p8_mult_21_n766, p8_mult_21_n765,
         p8_mult_21_n764, p8_mult_21_n763, p8_mult_21_n762, p8_mult_21_n761,
         p8_mult_21_n760, p8_mult_21_n759, p8_mult_21_n758, p8_mult_21_n756,
         p8_mult_21_n755, p8_mult_21_n754, p8_mult_21_n753, p8_mult_21_n752,
         p8_mult_21_n751, p8_mult_21_n750, p8_mult_21_n749, p8_mult_21_n748,
         p8_mult_21_n747, p8_mult_21_n746, p8_mult_21_n745, p8_mult_21_n744,
         p8_mult_21_n743, p8_mult_21_n742, p8_mult_21_n741, p8_mult_21_n739,
         p8_mult_21_n738, p8_mult_21_n737, p8_mult_21_n736, p8_mult_21_n735,
         p8_mult_21_n734, p8_mult_21_n733, p8_mult_21_n732, p8_mult_21_n731,
         p8_mult_21_n730, p8_mult_21_n729, p8_mult_21_n728, p8_mult_21_n727,
         p8_mult_21_n726, p8_mult_21_n725, p8_mult_21_n724, p8_mult_21_n722,
         p8_mult_21_n721, p8_mult_21_n720, p8_mult_21_n719, p8_mult_21_n718,
         p8_mult_21_n717, p8_mult_21_n716, p8_mult_21_n715, p8_mult_21_n714,
         p8_mult_21_n713, p8_mult_21_n712, p8_mult_21_n711, p8_mult_21_n710,
         p8_mult_21_n709, p8_mult_21_n708, p8_mult_21_n707, p8_mult_21_n706,
         p8_mult_21_n705, p8_mult_21_n704, p8_mult_21_n703, p8_mult_21_n702,
         p8_mult_21_n701, p8_mult_21_n700, p8_mult_21_n699, p8_mult_21_n698,
         p8_mult_21_n697, p8_mult_21_n696, p8_mult_21_n695, p8_mult_21_n694,
         p8_mult_21_n693, p8_mult_21_n692, p8_mult_21_n691, p8_mult_21_n690,
         p8_mult_21_n689, p8_mult_21_n688, p8_mult_21_n687, p8_mult_21_n686,
         p8_mult_21_n685, p8_mult_21_n682, p8_mult_21_n681, p8_mult_21_n670,
         p8_mult_21_n666, p8_mult_21_n657, p8_mult_21_n650, p8_mult_21_n646,
         p8_mult_21_n645, p8_mult_21_n644, p8_mult_21_n643, p8_mult_21_n641,
         p8_mult_21_n636, p8_mult_21_n419, p8_mult_21_n418, p8_mult_21_n417,
         p8_mult_21_n416, p8_mult_21_n415, p8_mult_21_n414, p8_mult_21_n413,
         p8_mult_21_n412, p8_mult_21_n411, p8_mult_21_n410, p8_mult_21_n409,
         p8_mult_21_n408, p8_mult_21_n406, p8_mult_21_n405, p8_mult_21_n404,
         p8_mult_21_n403, p8_mult_21_n402, p8_mult_21_n401, p8_mult_21_n400,
         p8_mult_21_n399, p8_mult_21_n398, p8_mult_21_n397, p8_mult_21_n396,
         p8_mult_21_n395, p8_mult_21_n394, p8_mult_21_n393, p8_mult_21_n390,
         p8_mult_21_n389, p8_mult_21_n388, p8_mult_21_n387, p8_mult_21_n386,
         p8_mult_21_n385, p8_mult_21_n384, p8_mult_21_n382, p8_mult_21_n381,
         p8_mult_21_n380, p8_mult_21_n379, p8_mult_21_n377, p8_mult_21_n376,
         p8_mult_21_n375, p8_mult_21_n374, p8_mult_21_n373, p8_mult_21_n372,
         p8_mult_21_n371, p8_mult_21_n370, p8_mult_21_n369, p8_mult_21_n368,
         p8_mult_21_n367, p8_mult_21_n366, p8_mult_21_n365, p8_mult_21_n363,
         p8_mult_21_n362, p8_mult_21_n361, p8_mult_21_n360, p8_mult_21_n359,
         p8_mult_21_n358, p8_mult_21_n357, p8_mult_21_n356, p8_mult_21_n355,
         p8_mult_21_n354, p8_mult_21_n353, p8_mult_21_n352, p8_mult_21_n351,
         p8_mult_21_n349, p8_mult_21_n348, p8_mult_21_n346, p8_mult_21_n345,
         p8_mult_21_n344, p8_mult_21_n343, p8_mult_21_n342, p8_mult_21_n341,
         p8_mult_21_n340, p8_mult_21_n339, p8_mult_21_n338, p8_mult_21_n337,
         p8_mult_21_n336, p8_mult_21_n335, p8_mult_21_n334, p8_mult_21_n333,
         p8_mult_21_n332, p8_mult_21_n331, p8_mult_21_n330, p8_mult_21_n329,
         p8_mult_21_n328, p8_mult_21_n327, p8_mult_21_n326, p8_mult_21_n325,
         p8_mult_21_n317, p8_mult_21_n316, p8_mult_21_n315, p8_mult_21_n314,
         p8_mult_21_n313, p8_mult_21_n312, p8_mult_21_n311, p8_mult_21_n308,
         p8_mult_21_n307, p8_mult_21_n304, p8_mult_21_n303, p8_mult_21_n302,
         p8_mult_21_n301, p8_mult_21_n300, p8_mult_21_n299, p8_mult_21_n298,
         p8_mult_21_n297, p8_mult_21_n296, p8_mult_21_n295, p8_mult_21_n294,
         p8_mult_21_n293, p8_mult_21_n292, p8_mult_21_n291, p8_mult_21_n290,
         p8_mult_21_n289, p8_mult_21_n284, p8_mult_21_n283, p8_mult_21_n282,
         p8_mult_21_n281, p8_mult_21_n280, p8_mult_21_n279, p8_mult_21_n276,
         p8_mult_21_n275, p8_mult_21_n274, p8_mult_21_n273, p8_mult_21_n272,
         p8_mult_21_n271, p8_mult_21_n270, p8_mult_21_n269, p8_mult_21_n268,
         p8_mult_21_n267, p8_mult_21_n266, p8_mult_21_n265, p8_mult_21_n264,
         p8_mult_21_n263, p8_mult_21_n262, p8_mult_21_n261, p8_mult_21_n260,
         p8_mult_21_n259, p8_mult_21_n258, p8_mult_21_n257, p8_mult_21_n256,
         p8_mult_21_n255, p8_mult_21_n254, p8_mult_21_n253, p8_mult_21_n252,
         p8_mult_21_n251, p8_mult_21_n250, p8_mult_21_n249, p8_mult_21_n248,
         p8_mult_21_n247, p8_mult_21_n246, p8_mult_21_n245, p8_mult_21_n244,
         p8_mult_21_n243, p8_mult_21_n242, p8_mult_21_n241, p8_mult_21_n240,
         p8_mult_21_n239, p8_mult_21_n238, p8_mult_21_n237, p8_mult_21_n236,
         p8_mult_21_n235, p8_mult_21_n234, p8_mult_21_n233, p8_mult_21_n232,
         p8_mult_21_n231, p8_mult_21_n230, p8_mult_21_n229, p8_mult_21_n228,
         p8_mult_21_n227, p8_mult_21_n226, p8_mult_21_n225, p8_mult_21_n224,
         p8_mult_21_n223, p8_mult_21_n222, p8_mult_21_n221, p8_mult_21_n220,
         p8_mult_21_n219, p8_mult_21_n218, p8_mult_21_n217, p8_mult_21_n216,
         p8_mult_21_n215, p8_mult_21_n214, p8_mult_21_n213, p8_mult_21_n212,
         p8_mult_21_n211, p8_mult_21_n210, p8_mult_21_n209, p8_mult_21_n208,
         p8_mult_21_n207, p8_mult_21_n206, p8_mult_21_n205, p8_mult_21_n204,
         p8_mult_21_n203, p8_mult_21_n202, p8_mult_21_n201, p8_mult_21_n200,
         p8_mult_21_n199, p8_mult_21_n198, p8_mult_21_n197, p8_mult_21_n196,
         p8_mult_21_n195, p8_mult_21_n194, p8_mult_21_n193, p8_mult_21_n192,
         p8_mult_21_n191, p8_mult_21_n190, p8_mult_21_n189, p8_mult_21_n188,
         p8_mult_21_n187, p8_mult_21_n186, p8_mult_21_n185, p8_mult_21_n184,
         p8_mult_21_n183, p8_mult_21_n182, p8_mult_21_n181, p8_mult_21_n180,
         p8_mult_21_n179, p8_mult_21_n178, p8_mult_21_n177, p8_mult_21_n176,
         p8_mult_21_n175, p8_mult_21_n174, p8_mult_21_n173, p8_mult_21_n172,
         p8_mult_21_n171, p8_mult_21_n170, p8_mult_21_n169, p8_mult_21_n168,
         p8_mult_21_n167, p8_mult_21_n166, p8_mult_21_n165, p8_mult_21_n164,
         p8_mult_21_n163, p8_mult_21_n162, p8_mult_21_n148, p8_mult_21_n147,
         p8_mult_21_n146, p8_mult_21_n145, p8_mult_21_n144, p8_mult_21_n143,
         p8_mult_21_n142, p8_mult_21_n141, p8_mult_21_n140, p8_mult_21_n139,
         p8_mult_21_n138, p8_mult_21_n137, p8_mult_21_n136, p9_mult_21_n927,
         p9_mult_21_n968, p9_mult_21_n1397, p9_mult_21_n1396, p9_mult_21_n1395,
         p9_mult_21_n1394, p9_mult_21_n1393, p9_mult_21_n1392,
         p9_mult_21_n1391, p9_mult_21_n1390, p9_mult_21_n1389,
         p9_mult_21_n1388, p9_mult_21_n1387, p9_mult_21_n1386,
         p9_mult_21_n1385, p9_mult_21_n1384, p9_mult_21_n1383,
         p9_mult_21_n1382, p9_mult_21_n1381, p9_mult_21_n1380,
         p9_mult_21_n1379, p9_mult_21_n1378, p9_mult_21_n1377,
         p9_mult_21_n1376, p9_mult_21_n1375, p9_mult_21_n1374,
         p9_mult_21_n1373, p9_mult_21_n1372, p9_mult_21_n1371,
         p9_mult_21_n1370, p9_mult_21_n1369, p9_mult_21_n1368,
         p9_mult_21_n1367, p9_mult_21_n1366, p9_mult_21_n1365,
         p9_mult_21_n1364, p9_mult_21_n1363, p9_mult_21_n1362,
         p9_mult_21_n1361, p9_mult_21_n1360, p9_mult_21_n1359,
         p9_mult_21_n1358, p9_mult_21_n1357, p9_mult_21_n1356,
         p9_mult_21_n1355, p9_mult_21_n1354, p9_mult_21_n1353,
         p9_mult_21_n1352, p9_mult_21_n1351, p9_mult_21_n1350,
         p9_mult_21_n1349, p9_mult_21_n1348, p9_mult_21_n1347,
         p9_mult_21_n1346, p9_mult_21_n1345, p9_mult_21_n1344,
         p9_mult_21_n1343, p9_mult_21_n1342, p9_mult_21_n1341,
         p9_mult_21_n1340, p9_mult_21_n1339, p9_mult_21_n1338,
         p9_mult_21_n1337, p9_mult_21_n1336, p9_mult_21_n1335,
         p9_mult_21_n1334, p9_mult_21_n1333, p9_mult_21_n1332,
         p9_mult_21_n1331, p9_mult_21_n1330, p9_mult_21_n1329,
         p9_mult_21_n1328, p9_mult_21_n1327, p9_mult_21_n1326,
         p9_mult_21_n1325, p9_mult_21_n1324, p9_mult_21_n1323,
         p9_mult_21_n1322, p9_mult_21_n1321, p9_mult_21_n1318,
         p9_mult_21_n1317, p9_mult_21_n1316, p9_mult_21_n1315,
         p9_mult_21_n1314, p9_mult_21_n1313, p9_mult_21_n1312,
         p9_mult_21_n1311, p9_mult_21_n1309, p9_mult_21_n1308,
         p9_mult_21_n1307, p9_mult_21_n1305, p9_mult_21_n1304,
         p9_mult_21_n1303, p9_mult_21_n1302, p9_mult_21_n1301,
         p9_mult_21_n1300, p9_mult_21_n1299, p9_mult_21_n1297,
         p9_mult_21_n1296, p9_mult_21_n1295, p9_mult_21_n1294,
         p9_mult_21_n1293, p9_mult_21_n1292, p9_mult_21_n1291,
         p9_mult_21_n1290, p9_mult_21_n1289, p9_mult_21_n1288,
         p9_mult_21_n1286, p9_mult_21_n1285, p9_mult_21_n1284,
         p9_mult_21_n1283, p9_mult_21_n1282, p9_mult_21_n1281,
         p9_mult_21_n1280, p9_mult_21_n1279, p9_mult_21_n1278,
         p9_mult_21_n1277, p9_mult_21_n1276, p9_mult_21_n1275,
         p9_mult_21_n1274, p9_mult_21_n1273, p9_mult_21_n1272,
         p9_mult_21_n1271, p9_mult_21_n1270, p9_mult_21_n1269,
         p9_mult_21_n1268, p9_mult_21_n1267, p9_mult_21_n1266,
         p9_mult_21_n1265, p9_mult_21_n1264, p9_mult_21_n1263,
         p9_mult_21_n1262, p9_mult_21_n1261, p9_mult_21_n1260,
         p9_mult_21_n1259, p9_mult_21_n1258, p9_mult_21_n1257,
         p9_mult_21_n1256, p9_mult_21_n1255, p9_mult_21_n1254,
         p9_mult_21_n1253, p9_mult_21_n1252, p9_mult_21_n1251,
         p9_mult_21_n1250, p9_mult_21_n1249, p9_mult_21_n1248,
         p9_mult_21_n1247, p9_mult_21_n1246, p9_mult_21_n1245,
         p9_mult_21_n1244, p9_mult_21_n1242, p9_mult_21_n1241,
         p9_mult_21_n1240, p9_mult_21_n1239, p9_mult_21_n1238,
         p9_mult_21_n1237, p9_mult_21_n1236, p9_mult_21_n1235,
         p9_mult_21_n1234, p9_mult_21_n1233, p9_mult_21_n1232,
         p9_mult_21_n1231, p9_mult_21_n1230, p9_mult_21_n1229,
         p9_mult_21_n1228, p9_mult_21_n1227, p9_mult_21_n1226,
         p9_mult_21_n1225, p9_mult_21_n1224, p9_mult_21_n1223,
         p9_mult_21_n1222, p9_mult_21_n1221, p9_mult_21_n1220,
         p9_mult_21_n1219, p9_mult_21_n1218, p9_mult_21_n1217,
         p9_mult_21_n1216, p9_mult_21_n1215, p9_mult_21_n1214,
         p9_mult_21_n1213, p9_mult_21_n1212, p9_mult_21_n1211,
         p9_mult_21_n1210, p9_mult_21_n1209, p9_mult_21_n1208,
         p9_mult_21_n1207, p9_mult_21_n1206, p9_mult_21_n1205,
         p9_mult_21_n1204, p9_mult_21_n1203, p9_mult_21_n1202,
         p9_mult_21_n1201, p9_mult_21_n1200, p9_mult_21_n1199,
         p9_mult_21_n1198, p9_mult_21_n1197, p9_mult_21_n1196,
         p9_mult_21_n1195, p9_mult_21_n1194, p9_mult_21_n1193,
         p9_mult_21_n1192, p9_mult_21_n1191, p9_mult_21_n1190,
         p9_mult_21_n1189, p9_mult_21_n1188, p9_mult_21_n1187,
         p9_mult_21_n1186, p9_mult_21_n1185, p9_mult_21_n1184,
         p9_mult_21_n1183, p9_mult_21_n1182, p9_mult_21_n1181,
         p9_mult_21_n1180, p9_mult_21_n1179, p9_mult_21_n1178,
         p9_mult_21_n1177, p9_mult_21_n1176, p9_mult_21_n1175,
         p9_mult_21_n1174, p9_mult_21_n1173, p9_mult_21_n1172,
         p9_mult_21_n1171, p9_mult_21_n1170, p9_mult_21_n1169,
         p9_mult_21_n1168, p9_mult_21_n1167, p9_mult_21_n1166,
         p9_mult_21_n1165, p9_mult_21_n1164, p9_mult_21_n1163,
         p9_mult_21_n1162, p9_mult_21_n1161, p9_mult_21_n1160,
         p9_mult_21_n1159, p9_mult_21_n1158, p9_mult_21_n1157,
         p9_mult_21_n1156, p9_mult_21_n1155, p9_mult_21_n1154,
         p9_mult_21_n1153, p9_mult_21_n1152, p9_mult_21_n1151,
         p9_mult_21_n1150, p9_mult_21_n1149, p9_mult_21_n1148,
         p9_mult_21_n1147, p9_mult_21_n1146, p9_mult_21_n1145,
         p9_mult_21_n1144, p9_mult_21_n1143, p9_mult_21_n1142,
         p9_mult_21_n1140, p9_mult_21_n1139, p9_mult_21_n1138,
         p9_mult_21_n1137, p9_mult_21_n1136, p9_mult_21_n1135,
         p9_mult_21_n1134, p9_mult_21_n1133, p9_mult_21_n1132,
         p9_mult_21_n1131, p9_mult_21_n1130, p9_mult_21_n1129,
         p9_mult_21_n1128, p9_mult_21_n1127, p9_mult_21_n1126,
         p9_mult_21_n1125, p9_mult_21_n1124, p9_mult_21_n1123,
         p9_mult_21_n1122, p9_mult_21_n1121, p9_mult_21_n1120,
         p9_mult_21_n1119, p9_mult_21_n1118, p9_mult_21_n1117,
         p9_mult_21_n1116, p9_mult_21_n1115, p9_mult_21_n1114,
         p9_mult_21_n1113, p9_mult_21_n1112, p9_mult_21_n1111,
         p9_mult_21_n1110, p9_mult_21_n1109, p9_mult_21_n1108,
         p9_mult_21_n1107, p9_mult_21_n1106, p9_mult_21_n1105,
         p9_mult_21_n1104, p9_mult_21_n1103, p9_mult_21_n1102,
         p9_mult_21_n1101, p9_mult_21_n1100, p9_mult_21_n1099,
         p9_mult_21_n1098, p9_mult_21_n1097, p9_mult_21_n1096,
         p9_mult_21_n1095, p9_mult_21_n1094, p9_mult_21_n1093,
         p9_mult_21_n1092, p9_mult_21_n1091, p9_mult_21_n1090,
         p9_mult_21_n1089, p9_mult_21_n1088, p9_mult_21_n1087,
         p9_mult_21_n1086, p9_mult_21_n1085, p9_mult_21_n1084,
         p9_mult_21_n1083, p9_mult_21_n1082, p9_mult_21_n1081,
         p9_mult_21_n1080, p9_mult_21_n1079, p9_mult_21_n1078,
         p9_mult_21_n1077, p9_mult_21_n1076, p9_mult_21_n1075,
         p9_mult_21_n1074, p9_mult_21_n1073, p9_mult_21_n1072,
         p9_mult_21_n1071, p9_mult_21_n1070, p9_mult_21_n1069,
         p9_mult_21_n1068, p9_mult_21_n1067, p9_mult_21_n1066,
         p9_mult_21_n1065, p9_mult_21_n1064, p9_mult_21_n1063,
         p9_mult_21_n1062, p9_mult_21_n1061, p9_mult_21_n1060,
         p9_mult_21_n1059, p9_mult_21_n1058, p9_mult_21_n1057,
         p9_mult_21_n1056, p9_mult_21_n1055, p9_mult_21_n1054,
         p9_mult_21_n1053, p9_mult_21_n1052, p9_mult_21_n1051,
         p9_mult_21_n1050, p9_mult_21_n1049, p9_mult_21_n1048,
         p9_mult_21_n1047, p9_mult_21_n1046, p9_mult_21_n1045,
         p9_mult_21_n1044, p9_mult_21_n1043, p9_mult_21_n1042,
         p9_mult_21_n1041, p9_mult_21_n1040, p9_mult_21_n1039,
         p9_mult_21_n1038, p9_mult_21_n1037, p9_mult_21_n1036,
         p9_mult_21_n1035, p9_mult_21_n1034, p9_mult_21_n1033,
         p9_mult_21_n1032, p9_mult_21_n1031, p9_mult_21_n1030,
         p9_mult_21_n1029, p9_mult_21_n1028, p9_mult_21_n1027,
         p9_mult_21_n1026, p9_mult_21_n1025, p9_mult_21_n1024,
         p9_mult_21_n1023, p9_mult_21_n1022, p9_mult_21_n1021,
         p9_mult_21_n1020, p9_mult_21_n1019, p9_mult_21_n1018,
         p9_mult_21_n1017, p9_mult_21_n1016, p9_mult_21_n1015,
         p9_mult_21_n1014, p9_mult_21_n1013, p9_mult_21_n1012,
         p9_mult_21_n1011, p9_mult_21_n1010, p9_mult_21_n1009,
         p9_mult_21_n1008, p9_mult_21_n1007, p9_mult_21_n1006,
         p9_mult_21_n1005, p9_mult_21_n1004, p9_mult_21_n1003,
         p9_mult_21_n1002, p9_mult_21_n1001, p9_mult_21_n1000, p9_mult_21_n999,
         p9_mult_21_n998, p9_mult_21_n997, p9_mult_21_n996, p9_mult_21_n995,
         p9_mult_21_n994, p9_mult_21_n993, p9_mult_21_n992, p9_mult_21_n991,
         p9_mult_21_n990, p9_mult_21_n989, p9_mult_21_n988, p9_mult_21_n987,
         p9_mult_21_n986, p9_mult_21_n985, p9_mult_21_n984, p9_mult_21_n983,
         p9_mult_21_n982, p9_mult_21_n981, p9_mult_21_n980, p9_mult_21_n979,
         p9_mult_21_n978, p9_mult_21_n977, p9_mult_21_n976, p9_mult_21_n975,
         p9_mult_21_n974, p9_mult_21_n973, p9_mult_21_n972, p9_mult_21_n971,
         p9_mult_21_n970, p9_mult_21_n969, p9_mult_21_n967, p9_mult_21_n966,
         p9_mult_21_n965, p9_mult_21_n964, p9_mult_21_n963, p9_mult_21_n962,
         p9_mult_21_n961, p9_mult_21_n960, p9_mult_21_n959, p9_mult_21_n958,
         p9_mult_21_n957, p9_mult_21_n956, p9_mult_21_n955, p9_mult_21_n954,
         p9_mult_21_n953, p9_mult_21_n952, p9_mult_21_n951, p9_mult_21_n950,
         p9_mult_21_n949, p9_mult_21_n948, p9_mult_21_n947, p9_mult_21_n946,
         p9_mult_21_n945, p9_mult_21_n944, p9_mult_21_n943, p9_mult_21_n942,
         p9_mult_21_n941, p9_mult_21_n940, p9_mult_21_n939, p9_mult_21_n938,
         p9_mult_21_n937, p9_mult_21_n936, p9_mult_21_n935, p9_mult_21_n934,
         p9_mult_21_n933, p9_mult_21_n932, p9_mult_21_n931, p9_mult_21_n930,
         p9_mult_21_n929, p9_mult_21_n928, p9_mult_21_n926, p9_mult_21_n925,
         p9_mult_21_n924, p9_mult_21_n923, p9_mult_21_n922, p9_mult_21_n921,
         p9_mult_21_n920, p9_mult_21_n919, p9_mult_21_n918, p9_mult_21_n917,
         p9_mult_21_n916, p9_mult_21_n915, p9_mult_21_n914, p9_mult_21_n913,
         p9_mult_21_n912, p9_mult_21_n911, p9_mult_21_n910, p9_mult_21_n909,
         p9_mult_21_n908, p9_mult_21_n907, p9_mult_21_n906, p9_mult_21_n905,
         p9_mult_21_n904, p9_mult_21_n903, p9_mult_21_n902, p9_mult_21_n901,
         p9_mult_21_n900, p9_mult_21_n899, p9_mult_21_n898, p9_mult_21_n897,
         p9_mult_21_n896, p9_mult_21_n895, p9_mult_21_n894, p9_mult_21_n893,
         p9_mult_21_n892, p9_mult_21_n890, p9_mult_21_n889, p9_mult_21_n888,
         p9_mult_21_n887, p9_mult_21_n886, p9_mult_21_n885, p9_mult_21_n883,
         p9_mult_21_n882, p9_mult_21_n881, p9_mult_21_n880, p9_mult_21_n879,
         p9_mult_21_n878, p9_mult_21_n877, p9_mult_21_n876, p9_mult_21_n875,
         p9_mult_21_n874, p9_mult_21_n873, p9_mult_21_n872, p9_mult_21_n871,
         p9_mult_21_n870, p9_mult_21_n869, p9_mult_21_n868, p9_mult_21_n867,
         p9_mult_21_n866, p9_mult_21_n865, p9_mult_21_n864, p9_mult_21_n863,
         p9_mult_21_n862, p9_mult_21_n860, p9_mult_21_n857, p9_mult_21_n845,
         p9_mult_21_n844, p9_mult_21_n843, p9_mult_21_n842, p9_mult_21_n841,
         p9_mult_21_n840, p9_mult_21_n839, p9_mult_21_n838, p11_mult_21_n845,
         p11_mult_21_n844, p11_mult_21_n843, p11_mult_21_n842,
         p11_mult_21_n841, p11_mult_21_n840, p11_mult_21_n839,
         p11_mult_21_n838, p11_mult_21_n832, p11_mult_21_n831,
         p11_mult_21_n830, p11_mult_21_n829, p11_mult_21_n828,
         p11_mult_21_n827, p11_mult_21_n826, p11_mult_21_n825,
         p11_mult_21_n824, p11_mult_21_n823, p11_mult_21_n822,
         p11_mult_21_n820, p11_mult_21_n819, p11_mult_21_n818,
         p11_mult_21_n817, p11_mult_21_n811, p11_mult_21_n807,
         p11_mult_21_n806, p11_mult_21_n805, p11_mult_21_n804,
         p11_mult_21_n803, p11_mult_21_n802, p11_mult_21_n801,
         p11_mult_21_n800, p11_mult_21_n799, p11_mult_21_n798,
         p11_mult_21_n797, p11_mult_21_n796, p11_mult_21_n795,
         p11_mult_21_n794, p11_mult_21_n793, p11_mult_21_n792,
         p11_mult_21_n791, p11_mult_21_n790, p11_mult_21_n789,
         p11_mult_21_n788, p11_mult_21_n787, p11_mult_21_n786,
         p11_mult_21_n785, p11_mult_21_n784, p11_mult_21_n783,
         p11_mult_21_n782, p11_mult_21_n781, p11_mult_21_n780,
         p11_mult_21_n779, p11_mult_21_n778, p11_mult_21_n777,
         p11_mult_21_n775, p11_mult_21_n774, p11_mult_21_n773,
         p11_mult_21_n772, p11_mult_21_n771, p11_mult_21_n770,
         p11_mult_21_n769, p11_mult_21_n768, p11_mult_21_n767,
         p11_mult_21_n766, p11_mult_21_n765, p11_mult_21_n764,
         p11_mult_21_n763, p11_mult_21_n762, p11_mult_21_n761,
         p11_mult_21_n760, p11_mult_21_n758, p11_mult_21_n757,
         p11_mult_21_n756, p11_mult_21_n755, p11_mult_21_n754,
         p11_mult_21_n753, p11_mult_21_n752, p11_mult_21_n751,
         p11_mult_21_n750, p11_mult_21_n749, p11_mult_21_n748,
         p11_mult_21_n747, p11_mult_21_n746, p11_mult_21_n745,
         p11_mult_21_n744, p11_mult_21_n743, p11_mult_21_n742,
         p11_mult_21_n741, p11_mult_21_n740, p11_mult_21_n739,
         p11_mult_21_n738, p11_mult_21_n737, p11_mult_21_n736,
         p11_mult_21_n735, p11_mult_21_n734, p11_mult_21_n733,
         p11_mult_21_n732, p11_mult_21_n731, p11_mult_21_n730,
         p11_mult_21_n729, p11_mult_21_n728, p11_mult_21_n727,
         p11_mult_21_n726, p11_mult_21_n724, p11_mult_21_n723,
         p11_mult_21_n722, p11_mult_21_n721, p11_mult_21_n720,
         p11_mult_21_n719, p11_mult_21_n718, p11_mult_21_n717,
         p11_mult_21_n716, p11_mult_21_n715, p11_mult_21_n714,
         p11_mult_21_n713, p11_mult_21_n712, p11_mult_21_n711,
         p11_mult_21_n710, p11_mult_21_n709, p11_mult_21_n708,
         p11_mult_21_n707, p11_mult_21_n706, p11_mult_21_n704,
         p11_mult_21_n703, p11_mult_21_n702, p11_mult_21_n701,
         p11_mult_21_n700, p11_mult_21_n699, p11_mult_21_n698,
         p11_mult_21_n697, p11_mult_21_n696, p11_mult_21_n695,
         p11_mult_21_n694, p11_mult_21_n693, p11_mult_21_n692,
         p11_mult_21_n691, p11_mult_21_n690, p11_mult_21_n689,
         p11_mult_21_n688, p11_mult_21_n687, p11_mult_21_n682,
         p11_mult_21_n681, p11_mult_21_n680, p11_mult_21_n679,
         p11_mult_21_n672, p11_mult_21_n671, p11_mult_21_n670,
         p11_mult_21_n669, p11_mult_21_n668, p11_mult_21_n662,
         p11_mult_21_n661, p11_mult_21_n660, p11_mult_21_n659,
         p11_mult_21_n652, p11_mult_21_n651, p11_mult_21_n646,
         p11_mult_21_n642, p11_mult_21_n641, p11_mult_21_n640,
         p11_mult_21_n636, p11_mult_21_n635, p11_mult_21_n418,
         p11_mult_21_n417, p11_mult_21_n416, p11_mult_21_n415,
         p11_mult_21_n414, p11_mult_21_n413, p11_mult_21_n412,
         p11_mult_21_n411, p11_mult_21_n410, p11_mult_21_n409,
         p11_mult_21_n408, p11_mult_21_n405, p11_mult_21_n404,
         p11_mult_21_n403, p11_mult_21_n402, p11_mult_21_n401,
         p11_mult_21_n400, p11_mult_21_n399, p11_mult_21_n398,
         p11_mult_21_n397, p11_mult_21_n396, p11_mult_21_n395,
         p11_mult_21_n394, p11_mult_21_n393, p11_mult_21_n390,
         p11_mult_21_n389, p11_mult_21_n388, p11_mult_21_n387,
         p11_mult_21_n386, p11_mult_21_n385, p11_mult_21_n384,
         p11_mult_21_n382, p11_mult_21_n381, p11_mult_21_n380,
         p11_mult_21_n379, p11_mult_21_n378, p11_mult_21_n377,
         p11_mult_21_n376, p11_mult_21_n375, p11_mult_21_n374,
         p11_mult_21_n373, p11_mult_21_n372, p11_mult_21_n371,
         p11_mult_21_n370, p11_mult_21_n369, p11_mult_21_n368,
         p11_mult_21_n367, p11_mult_21_n366, p11_mult_21_n365,
         p11_mult_21_n363, p11_mult_21_n362, p11_mult_21_n361,
         p11_mult_21_n360, p11_mult_21_n359, p11_mult_21_n358,
         p11_mult_21_n357, p11_mult_21_n356, p11_mult_21_n355,
         p11_mult_21_n354, p11_mult_21_n353, p11_mult_21_n352,
         p11_mult_21_n351, p11_mult_21_n349, p11_mult_21_n348,
         p11_mult_21_n346, p11_mult_21_n345, p11_mult_21_n344,
         p11_mult_21_n343, p11_mult_21_n342, p11_mult_21_n341,
         p11_mult_21_n340, p11_mult_21_n339, p11_mult_21_n338,
         p11_mult_21_n337, p11_mult_21_n336, p11_mult_21_n335,
         p11_mult_21_n334, p11_mult_21_n333, p11_mult_21_n332,
         p11_mult_21_n331, p11_mult_21_n330, p11_mult_21_n329,
         p11_mult_21_n328, p11_mult_21_n327, p11_mult_21_n326,
         p11_mult_21_n325, p11_mult_21_n320, p11_mult_21_n317,
         p11_mult_21_n314, p11_mult_21_n313, p11_mult_21_n312,
         p11_mult_21_n311, p11_mult_21_n308, p11_mult_21_n307,
         p11_mult_21_n304, p11_mult_21_n303, p11_mult_21_n302,
         p11_mult_21_n301, p11_mult_21_n300, p11_mult_21_n299,
         p11_mult_21_n298, p11_mult_21_n297, p11_mult_21_n296,
         p11_mult_21_n295, p11_mult_21_n294, p11_mult_21_n293,
         p11_mult_21_n292, p11_mult_21_n291, p11_mult_21_n290,
         p11_mult_21_n289, p11_mult_21_n288, p11_mult_21_n287,
         p11_mult_21_n286, p11_mult_21_n285, p11_mult_21_n284,
         p11_mult_21_n283, p11_mult_21_n282, p11_mult_21_n281,
         p11_mult_21_n280, p11_mult_21_n279, p11_mult_21_n278,
         p11_mult_21_n277, p11_mult_21_n276, p11_mult_21_n275,
         p11_mult_21_n274, p11_mult_21_n273, p11_mult_21_n272,
         p11_mult_21_n271, p11_mult_21_n270, p11_mult_21_n269,
         p11_mult_21_n268, p11_mult_21_n267, p11_mult_21_n266,
         p11_mult_21_n265, p11_mult_21_n264, p11_mult_21_n263,
         p11_mult_21_n262, p11_mult_21_n261, p11_mult_21_n260,
         p11_mult_21_n259, p11_mult_21_n258, p11_mult_21_n257,
         p11_mult_21_n256, p11_mult_21_n255, p11_mult_21_n254,
         p11_mult_21_n253, p11_mult_21_n252, p11_mult_21_n251,
         p11_mult_21_n250, p11_mult_21_n249, p11_mult_21_n248,
         p11_mult_21_n247, p11_mult_21_n246, p11_mult_21_n245,
         p11_mult_21_n244, p11_mult_21_n243, p11_mult_21_n242,
         p11_mult_21_n241, p11_mult_21_n240, p11_mult_21_n239,
         p11_mult_21_n238, p11_mult_21_n237, p11_mult_21_n236,
         p11_mult_21_n235, p11_mult_21_n234, p11_mult_21_n233,
         p11_mult_21_n232, p11_mult_21_n231, p11_mult_21_n230,
         p11_mult_21_n229, p11_mult_21_n228, p11_mult_21_n227,
         p11_mult_21_n226, p11_mult_21_n225, p11_mult_21_n224,
         p11_mult_21_n223, p11_mult_21_n222, p11_mult_21_n221,
         p11_mult_21_n220, p11_mult_21_n219, p11_mult_21_n218,
         p11_mult_21_n217, p11_mult_21_n216, p11_mult_21_n215,
         p11_mult_21_n214, p11_mult_21_n213, p11_mult_21_n212,
         p11_mult_21_n211, p11_mult_21_n210, p11_mult_21_n209,
         p11_mult_21_n208, p11_mult_21_n207, p11_mult_21_n206,
         p11_mult_21_n205, p11_mult_21_n204, p11_mult_21_n203,
         p11_mult_21_n202, p11_mult_21_n201, p11_mult_21_n200,
         p11_mult_21_n199, p11_mult_21_n198, p11_mult_21_n197,
         p11_mult_21_n196, p11_mult_21_n195, p11_mult_21_n194,
         p11_mult_21_n193, p11_mult_21_n192, p11_mult_21_n191,
         p11_mult_21_n190, p11_mult_21_n189, p11_mult_21_n188,
         p11_mult_21_n187, p11_mult_21_n186, p11_mult_21_n185,
         p11_mult_21_n184, p11_mult_21_n183, p11_mult_21_n182,
         p11_mult_21_n181, p11_mult_21_n180, p11_mult_21_n179,
         p11_mult_21_n178, p11_mult_21_n177, p11_mult_21_n176,
         p11_mult_21_n175, p11_mult_21_n174, p11_mult_21_n173,
         p11_mult_21_n172, p11_mult_21_n171, p11_mult_21_n170,
         p11_mult_21_n169, p11_mult_21_n168, p11_mult_21_n167,
         p11_mult_21_n166, p11_mult_21_n165, p11_mult_21_n164,
         p11_mult_21_n163, p11_mult_21_n162, p11_mult_21_n148,
         p11_mult_21_n146, p11_mult_21_n145, p11_mult_21_n144,
         p11_mult_21_n143, p11_mult_21_n142, p11_mult_21_n141,
         p11_mult_21_n140, p11_mult_21_n139, p11_mult_21_n138,
         p11_mult_21_n137, p11_mult_21_n136, p10_mult_21_n968,
         p10_mult_21_n1396, p10_mult_21_n1392, p10_mult_21_n1391,
         p10_mult_21_n1390, p10_mult_21_n1389, p10_mult_21_n1388,
         p10_mult_21_n1387, p10_mult_21_n1386, p10_mult_21_n1385,
         p10_mult_21_n1384, p10_mult_21_n1383, p10_mult_21_n1382,
         p10_mult_21_n1381, p10_mult_21_n1380, p10_mult_21_n1378,
         p10_mult_21_n1377, p10_mult_21_n1376, p10_mult_21_n1375,
         p10_mult_21_n1374, p10_mult_21_n1373, p10_mult_21_n1372,
         p10_mult_21_n1371, p10_mult_21_n1369, p10_mult_21_n1368,
         p10_mult_21_n1367, p10_mult_21_n1366, p10_mult_21_n1365,
         p10_mult_21_n1364, p10_mult_21_n1363, p10_mult_21_n1362,
         p10_mult_21_n1361, p10_mult_21_n1360, p10_mult_21_n1359,
         p10_mult_21_n1358, p10_mult_21_n1357, p10_mult_21_n1356,
         p10_mult_21_n1355, p10_mult_21_n1354, p10_mult_21_n1353,
         p10_mult_21_n1352, p10_mult_21_n1351, p10_mult_21_n1350,
         p10_mult_21_n1349, p10_mult_21_n1348, p10_mult_21_n1347,
         p10_mult_21_n1346, p10_mult_21_n1345, p10_mult_21_n1344,
         p10_mult_21_n1343, p10_mult_21_n1342, p10_mult_21_n1341,
         p10_mult_21_n1340, p10_mult_21_n1337, p10_mult_21_n1336,
         p10_mult_21_n1335, p10_mult_21_n1334, p10_mult_21_n1333,
         p10_mult_21_n1332, p10_mult_21_n1331, p10_mult_21_n1330,
         p10_mult_21_n1329, p10_mult_21_n1328, p10_mult_21_n1327,
         p10_mult_21_n1326, p10_mult_21_n1325, p10_mult_21_n1324,
         p10_mult_21_n1323, p10_mult_21_n1322, p10_mult_21_n1321,
         p10_mult_21_n1318, p10_mult_21_n1317, p10_mult_21_n1316,
         p10_mult_21_n1315, p10_mult_21_n1314, p10_mult_21_n1313,
         p10_mult_21_n1312, p10_mult_21_n1311, p10_mult_21_n1310,
         p10_mult_21_n1309, p10_mult_21_n1308, p10_mult_21_n1307,
         p10_mult_21_n1305, p10_mult_21_n1304, p10_mult_21_n1303,
         p10_mult_21_n1302, p10_mult_21_n1301, p10_mult_21_n1300,
         p10_mult_21_n1299, p10_mult_21_n1298, p10_mult_21_n1297,
         p10_mult_21_n1296, p10_mult_21_n1295, p10_mult_21_n1294,
         p10_mult_21_n1293, p10_mult_21_n1292, p10_mult_21_n1288,
         p10_mult_21_n1287, p10_mult_21_n1286, p10_mult_21_n1285,
         p10_mult_21_n1284, p10_mult_21_n1283, p10_mult_21_n1282,
         p10_mult_21_n1281, p10_mult_21_n1280, p10_mult_21_n1279,
         p10_mult_21_n1278, p10_mult_21_n1277, p10_mult_21_n1276,
         p10_mult_21_n1275, p10_mult_21_n1274, p10_mult_21_n1273,
         p10_mult_21_n1272, p10_mult_21_n1271, p10_mult_21_n1270,
         p10_mult_21_n1269, p10_mult_21_n1268, p10_mult_21_n1267,
         p10_mult_21_n1266, p10_mult_21_n1265, p10_mult_21_n1264,
         p10_mult_21_n1261, p10_mult_21_n1260, p10_mult_21_n1259,
         p10_mult_21_n1258, p10_mult_21_n1257, p10_mult_21_n1256,
         p10_mult_21_n1255, p10_mult_21_n1254, p10_mult_21_n1253,
         p10_mult_21_n1252, p10_mult_21_n1251, p10_mult_21_n1250,
         p10_mult_21_n1249, p10_mult_21_n1248, p10_mult_21_n1247,
         p10_mult_21_n1246, p10_mult_21_n1243, p10_mult_21_n1242,
         p10_mult_21_n1241, p10_mult_21_n1240, p10_mult_21_n1238,
         p10_mult_21_n1237, p10_mult_21_n1236, p10_mult_21_n1235,
         p10_mult_21_n1234, p10_mult_21_n1233, p10_mult_21_n1232,
         p10_mult_21_n1231, p10_mult_21_n1230, p10_mult_21_n1229,
         p10_mult_21_n1228, p10_mult_21_n1227, p10_mult_21_n1226,
         p10_mult_21_n1225, p10_mult_21_n1224, p10_mult_21_n1222,
         p10_mult_21_n1221, p10_mult_21_n1220, p10_mult_21_n1219,
         p10_mult_21_n1218, p10_mult_21_n1217, p10_mult_21_n1216,
         p10_mult_21_n1215, p10_mult_21_n1214, p10_mult_21_n1213,
         p10_mult_21_n1212, p10_mult_21_n1211, p10_mult_21_n1210,
         p10_mult_21_n1209, p10_mult_21_n1208, p10_mult_21_n1207,
         p10_mult_21_n1206, p10_mult_21_n1205, p10_mult_21_n1204,
         p10_mult_21_n1203, p10_mult_21_n1202, p10_mult_21_n1201,
         p10_mult_21_n1200, p10_mult_21_n1199, p10_mult_21_n1198,
         p10_mult_21_n1197, p10_mult_21_n1196, p10_mult_21_n1195,
         p10_mult_21_n1194, p10_mult_21_n1193, p10_mult_21_n1192,
         p10_mult_21_n1191, p10_mult_21_n1190, p10_mult_21_n1189,
         p10_mult_21_n1188, p10_mult_21_n1187, p10_mult_21_n1186,
         p10_mult_21_n1185, p10_mult_21_n1184, p10_mult_21_n1183,
         p10_mult_21_n1182, p10_mult_21_n1181, p10_mult_21_n1180,
         p10_mult_21_n1179, p10_mult_21_n1178, p10_mult_21_n1177,
         p10_mult_21_n1176, p10_mult_21_n1175, p10_mult_21_n1174,
         p10_mult_21_n1173, p10_mult_21_n1172, p10_mult_21_n1171,
         p10_mult_21_n1170, p10_mult_21_n1169, p10_mult_21_n1168,
         p10_mult_21_n1167, p10_mult_21_n1166, p10_mult_21_n1165,
         p10_mult_21_n1164, p10_mult_21_n1163, p10_mult_21_n1162,
         p10_mult_21_n1161, p10_mult_21_n1160, p10_mult_21_n1159,
         p10_mult_21_n1158, p10_mult_21_n1157, p10_mult_21_n1156,
         p10_mult_21_n1155, p10_mult_21_n1154, p10_mult_21_n1153,
         p10_mult_21_n1152, p10_mult_21_n1151, p10_mult_21_n1150,
         p10_mult_21_n1149, p10_mult_21_n1148, p10_mult_21_n1147,
         p10_mult_21_n1146, p10_mult_21_n1145, p10_mult_21_n1144,
         p10_mult_21_n1143, p10_mult_21_n1142, p10_mult_21_n1141,
         p10_mult_21_n1140, p10_mult_21_n1139, p10_mult_21_n1138,
         p10_mult_21_n1137, p10_mult_21_n1136, p10_mult_21_n1135,
         p10_mult_21_n1134, p10_mult_21_n1133, p10_mult_21_n1132,
         p10_mult_21_n1131, p10_mult_21_n1130, p10_mult_21_n1129,
         p10_mult_21_n1128, p10_mult_21_n1127, p10_mult_21_n1126,
         p10_mult_21_n1125, p10_mult_21_n1124, p10_mult_21_n1123,
         p10_mult_21_n1122, p10_mult_21_n1121, p10_mult_21_n1120,
         p10_mult_21_n1119, p10_mult_21_n1118, p10_mult_21_n1117,
         p10_mult_21_n1116, p10_mult_21_n1114, p10_mult_21_n1113,
         p10_mult_21_n1112, p10_mult_21_n1111, p10_mult_21_n1110,
         p10_mult_21_n1109, p10_mult_21_n1108, p10_mult_21_n1107,
         p10_mult_21_n1106, p10_mult_21_n1105, p10_mult_21_n1104,
         p10_mult_21_n1103, p10_mult_21_n1102, p10_mult_21_n1101,
         p10_mult_21_n1100, p10_mult_21_n1099, p10_mult_21_n1098,
         p10_mult_21_n1097, p10_mult_21_n1096, p10_mult_21_n1095,
         p10_mult_21_n1094, p10_mult_21_n1093, p10_mult_21_n1092,
         p10_mult_21_n1091, p10_mult_21_n1090, p10_mult_21_n1089,
         p10_mult_21_n1088, p10_mult_21_n1087, p10_mult_21_n1086,
         p10_mult_21_n1085, p10_mult_21_n1084, p10_mult_21_n1083,
         p10_mult_21_n1082, p10_mult_21_n1081, p10_mult_21_n1080,
         p10_mult_21_n1079, p10_mult_21_n1078, p10_mult_21_n1077,
         p10_mult_21_n1076, p10_mult_21_n1075, p10_mult_21_n1074,
         p10_mult_21_n1073, p10_mult_21_n1072, p10_mult_21_n1071,
         p10_mult_21_n1070, p10_mult_21_n1069, p10_mult_21_n1068,
         p10_mult_21_n1067, p10_mult_21_n1066, p10_mult_21_n1065,
         p10_mult_21_n1064, p10_mult_21_n1063, p10_mult_21_n1062,
         p10_mult_21_n1061, p10_mult_21_n1060, p10_mult_21_n1059,
         p10_mult_21_n1058, p10_mult_21_n1057, p10_mult_21_n1056,
         p10_mult_21_n1055, p10_mult_21_n1054, p10_mult_21_n1053,
         p10_mult_21_n1052, p10_mult_21_n1051, p10_mult_21_n1050,
         p10_mult_21_n1049, p10_mult_21_n1048, p10_mult_21_n1047,
         p10_mult_21_n1046, p10_mult_21_n1045, p10_mult_21_n1044,
         p10_mult_21_n1043, p10_mult_21_n1042, p10_mult_21_n1041,
         p10_mult_21_n1040, p10_mult_21_n1039, p10_mult_21_n1038,
         p10_mult_21_n1037, p10_mult_21_n1036, p10_mult_21_n1035,
         p10_mult_21_n1034, p10_mult_21_n1033, p10_mult_21_n1032,
         p10_mult_21_n1031, p10_mult_21_n1030, p10_mult_21_n1029,
         p10_mult_21_n1028, p10_mult_21_n1027, p10_mult_21_n1026,
         p10_mult_21_n1025, p10_mult_21_n1024, p10_mult_21_n1023,
         p10_mult_21_n1022, p10_mult_21_n1021, p10_mult_21_n1020,
         p10_mult_21_n1019, p10_mult_21_n1018, p10_mult_21_n1017,
         p10_mult_21_n1016, p10_mult_21_n1015, p10_mult_21_n1014,
         p10_mult_21_n1013, p10_mult_21_n1012, p10_mult_21_n1011,
         p10_mult_21_n1010, p10_mult_21_n1009, p10_mult_21_n1008,
         p10_mult_21_n1007, p10_mult_21_n1006, p10_mult_21_n1005,
         p10_mult_21_n1004, p10_mult_21_n1003, p10_mult_21_n1002,
         p10_mult_21_n1001, p10_mult_21_n1000, p10_mult_21_n999,
         p10_mult_21_n998, p10_mult_21_n997, p10_mult_21_n996,
         p10_mult_21_n995, p10_mult_21_n994, p10_mult_21_n993,
         p10_mult_21_n992, p10_mult_21_n991, p10_mult_21_n990,
         p10_mult_21_n989, p10_mult_21_n988, p10_mult_21_n986,
         p10_mult_21_n985, p10_mult_21_n984, p10_mult_21_n983,
         p10_mult_21_n982, p10_mult_21_n981, p10_mult_21_n980,
         p10_mult_21_n979, p10_mult_21_n978, p10_mult_21_n977,
         p10_mult_21_n976, p10_mult_21_n974, p10_mult_21_n973,
         p10_mult_21_n972, p10_mult_21_n971, p10_mult_21_n970,
         p10_mult_21_n969, p10_mult_21_n967, p10_mult_21_n966,
         p10_mult_21_n965, p10_mult_21_n964, p10_mult_21_n963,
         p10_mult_21_n962, p10_mult_21_n961, p10_mult_21_n960,
         p10_mult_21_n959, p10_mult_21_n958, p10_mult_21_n957,
         p10_mult_21_n956, p10_mult_21_n955, p10_mult_21_n954,
         p10_mult_21_n953, p10_mult_21_n952, p10_mult_21_n951,
         p10_mult_21_n950, p10_mult_21_n949, p10_mult_21_n948,
         p10_mult_21_n947, p10_mult_21_n946, p10_mult_21_n945,
         p10_mult_21_n944, p10_mult_21_n943, p10_mult_21_n942,
         p10_mult_21_n941, p10_mult_21_n940, p10_mult_21_n938,
         p10_mult_21_n937, p10_mult_21_n936, p10_mult_21_n935,
         p10_mult_21_n934, p10_mult_21_n933, p10_mult_21_n932,
         p10_mult_21_n931, p10_mult_21_n930, p10_mult_21_n929,
         p10_mult_21_n928, p10_mult_21_n927, p10_mult_21_n926,
         p10_mult_21_n925, p10_mult_21_n924, p10_mult_21_n923,
         p10_mult_21_n922, p10_mult_21_n921, p10_mult_21_n920,
         p10_mult_21_n919, p10_mult_21_n918, p10_mult_21_n917,
         p10_mult_21_n916, p10_mult_21_n915, p10_mult_21_n914,
         p10_mult_21_n913, p10_mult_21_n912, p10_mult_21_n911,
         p10_mult_21_n910, p10_mult_21_n909, p10_mult_21_n908,
         p10_mult_21_n907, p10_mult_21_n906, p10_mult_21_n904,
         p10_mult_21_n903, p10_mult_21_n902, p10_mult_21_n901,
         p10_mult_21_n900, p10_mult_21_n899, p10_mult_21_n898,
         p10_mult_21_n897, p10_mult_21_n896, p10_mult_21_n895,
         p10_mult_21_n894, p10_mult_21_n893, p10_mult_21_n892,
         p10_mult_21_n890, p10_mult_21_n889, p10_mult_21_n888,
         p10_mult_21_n887, p10_mult_21_n886, p10_mult_21_n885,
         p10_mult_21_n883, p10_mult_21_n882, p10_mult_21_n881,
         p10_mult_21_n880, p10_mult_21_n879, p10_mult_21_n878,
         p10_mult_21_n877, p10_mult_21_n875, p10_mult_21_n874,
         p10_mult_21_n873, p10_mult_21_n872, p10_mult_21_n871,
         p10_mult_21_n869, p10_mult_21_n868, p10_mult_21_n866,
         p10_mult_21_n864, p10_mult_21_n863, p10_mult_21_n862,
         p10_mult_21_n861, p10_mult_21_n860, p10_mult_21_n857,
         p10_mult_21_n849, p10_mult_21_n848, p10_mult_21_n845,
         p10_mult_21_n844, p10_mult_21_n843, p10_mult_21_n842,
         p10_mult_21_n841, p10_mult_21_n840, p10_mult_21_n839,
         p10_mult_21_n838, p10_mult_21_n837, p10_mult_21_n836,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_1_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_2_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_3_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_4_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_5_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_6_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_7_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_8_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_9_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_10_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_13_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_, s6_add_21_carry_1_,
         s6_add_21_carry_2_, s6_add_21_carry_3_, s6_add_21_carry_4_,
         s6_add_21_carry_5_, s6_add_21_carry_6_, s6_add_21_carry_7_,
         s6_add_21_carry_8_, s6_add_21_carry_9_, s6_add_21_carry_10_,
         s6_add_21_carry_11_, s6_add_21_carry_12_, s6_add_21_carry_13_,
         s7_add_21_carry_1_, s7_add_21_carry_2_, s7_add_21_carry_3_,
         s7_add_21_carry_4_, s7_add_21_carry_5_, s7_add_21_carry_6_,
         s7_add_21_carry_7_, s7_add_21_carry_8_, s7_add_21_carry_9_,
         s7_add_21_carry_10_, s7_add_21_carry_11_, s7_add_21_carry_12_,
         s7_add_21_carry_13_, s8_add_21_carry_1_, s8_add_21_carry_2_,
         s8_add_21_carry_3_, s8_add_21_carry_4_, s8_add_21_carry_5_,
         s8_add_21_carry_6_, s8_add_21_carry_7_, s8_add_21_carry_8_,
         s8_add_21_carry_9_, s8_add_21_carry_10_, s8_add_21_carry_11_,
         s8_add_21_carry_12_, s8_add_21_carry_13_, s9_add_21_carry_1_,
         s9_add_21_carry_2_, s9_add_21_carry_3_, s9_add_21_carry_4_,
         s9_add_21_carry_5_, s9_add_21_carry_6_, s9_add_21_carry_7_,
         s9_add_21_carry_8_, s9_add_21_carry_9_, s9_add_21_carry_10_,
         s9_add_21_carry_11_, s9_add_21_carry_12_, s9_add_21_carry_13_, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942;
  wire   [13:0] xin_in;
  wire   [13:0] xin;
  wire   [13:0] w;
  wire   [13:0] reg1_reg;
  wire   [13:0] temp1;
  wire   [13:0] mul1_reg;
  wire   [13:0] reg2;
  wire   [13:0] reg2_reg;
  wire   [13:0] temp2;
  wire   [13:0] mul2_reg;
  wire   [13:0] reg3;
  wire   [13:0] reg3_reg;
  wire   [13:0] temp3;
  wire   [13:0] mul3_reg;
  wire   [13:0] reg5;
  wire   [13:0] reg4_reg;
  wire   [13:0] temp4;
  wire   [13:0] mul4_reg;
  wire   [13:0] temp6;
  wire   [13:0] reg4;
  wire   [13:0] temp5;
  wire   [13:0] reg6;
  wire   [13:0] reg7;
  wire   [13:0] ff;

  reg_0 REGISTER_in ( .RST_n(RST_n), .VIN(VIN), .d({n66, n67, n68, n69, n70, 
        n74, n75, n76, n77, n78, n79, n71, n72, n73}), .CLK(CLK), .q(xin) );
  reg_7 REGISTER_out ( .RST_n(RST_n), .VIN(VIN), .d(ff), .CLK(CLK), .q(DOUT)
         );
  DFFR_X1 MY_CLK_r_REG0_S1 ( .D(n185), .CK(CLK), .RN(RST_n), .Q(VOUT), .QN(n30) );
  DFFR_X1 REG1_1_MY_CLK_r_REG3_S4 ( .D(REG1_1_n254), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[13]), .QN(n916) );
  DFFS_X1 REG2_1_MY_CLK_r_REG37_S16 ( .D(REG2_1_n272), .CK(CLK), .SN(RST_n), 
        .QN(REG2_1_n271) );
  DFFR_X1 REG2_1_MY_CLK_r_REG39_S15 ( .D(REG2_1_n259), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[11]), .QN(n917) );
  DFFS_X1 REG2_1_MY_CLK_r_REG36_S15 ( .D(REG2_1_n75), .CK(CLK), .SN(RST_n), 
        .QN(REG2_1_n92) );
  DFFR_X1 REG3_1_MY_CLK_r_REG53_S16 ( .D(REG3_1_n254), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[13]), .QN(n915) );
  DFFR_X1 REG4_1_MY_CLK_r_REG93_S20 ( .D(REG4_1_n254), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[12]), .QN(n918) );
  DFFS_X2 REG11_MY_CLK_r_REG123_S13 ( .D(REG11_n64), .CK(CLK), .SN(RST_n), .Q(
        n575), .QN(reg2[3]) );
  DFFR_X1 REG11_MY_CLK_r_REG113_S16 ( .D(REG11_n266), .CK(CLK), .RN(RST_n), 
        .Q(reg2[0]), .QN(p11_mult_21_n693) );
  DFFR_X1 REG11_MY_CLK_r_REG33_S13 ( .D(REG11_n263), .CK(CLK), .RN(RST_n), .Q(
        reg2[4]), .QN(n894) );
  DFFR_X1 REG11_MY_CLK_r_REG83_S16 ( .D(REG11_n264), .CK(CLK), .RN(RST_n), .Q(
        reg2[2]), .QN(n895) );
  DFFR_X1 REG11_MY_CLK_r_REG21_S5 ( .D(REG11_n255), .CK(CLK), .RN(RST_n), .Q(
        reg2[12]), .QN(n890) );
  DFFR_X1 REG11_MY_CLK_r_REG153_S11 ( .D(REG11_n261), .CK(CLK), .RN(RST_n), 
        .Q(reg2[6]), .QN(n893) );
  DFFR_X1 REG11_MY_CLK_r_REG27_S9 ( .D(REG11_n257), .CK(CLK), .RN(RST_n), .Q(
        reg2[10]), .QN(n891) );
  DFFR_X1 REG11_MY_CLK_r_REG137_S11 ( .D(REG11_n259), .CK(CLK), .RN(RST_n), 
        .Q(reg2[8]), .QN(n892) );
  DFFR_X1 REG21_MY_CLK_r_REG155_S12 ( .D(REG21_n260), .CK(CLK), .RN(RST_n), 
        .Q(reg3[6]), .QN(n927) );
  DFFR_X1 REG21_MY_CLK_r_REG163_S12 ( .D(REG21_n261), .CK(CLK), .RN(RST_n), 
        .Q(reg3[5]), .QN(n928) );
  DFFR_X1 REG21_MY_CLK_r_REG107_S17 ( .D(REG21_n265), .CK(CLK), .RN(RST_n), 
        .Q(reg3[1]), .QN(n931) );
  DFFR_X1 REG21_MY_CLK_r_REG51_S14 ( .D(REG21_n262), .CK(CLK), .RN(RST_n), .Q(
        reg3[4]), .QN(n929) );
  DFFR_X1 REG21_MY_CLK_r_REG85_S17 ( .D(REG21_n264), .CK(CLK), .RN(RST_n), .Q(
        reg3[2]), .QN(n930) );
  DFFR_X1 REG21_MY_CLK_r_REG125_S14 ( .D(REG21_n263), .CK(CLK), .RN(RST_n), 
        .Q(reg3[3]), .QN(n919) );
  DFFR_X1 REG21_MY_CLK_r_REG115_S17 ( .D(REG21_n266), .CK(CLK), .RN(RST_n), 
        .Q(reg3[0]), .QN(n932) );
  DFFR_X1 REG21_MY_CLK_r_REG194_S4 ( .D(REG21_n253), .CK(CLK), .RN(RST_n), .Q(
        reg3[13]), .QN(n920) );
  DFFR_X1 REG21_MY_CLK_r_REG182_S6 ( .D(REG21_n254), .CK(CLK), .RN(RST_n), .Q(
        reg3[12]), .QN(n921) );
  DFFR_X1 REG21_MY_CLK_r_REG176_S8 ( .D(REG21_n255), .CK(CLK), .RN(RST_n), .Q(
        reg3[11]), .QN(n922) );
  DFFR_X1 REG21_MY_CLK_r_REG169_S10 ( .D(REG21_n256), .CK(CLK), .RN(RST_n), 
        .Q(reg3[10]), .QN(n923) );
  DFFR_X1 REG21_MY_CLK_r_REG131_S12 ( .D(REG21_n257), .CK(CLK), .RN(RST_n), 
        .Q(reg3[9]), .QN(n924) );
  DFFR_X1 REG21_MY_CLK_r_REG139_S12 ( .D(REG21_n258), .CK(CLK), .RN(RST_n), 
        .Q(reg3[8]), .QN(n925) );
  DFFR_X1 REG21_MY_CLK_r_REG147_S12 ( .D(REG21_n259), .CK(CLK), .RN(RST_n), 
        .Q(reg3[7]), .QN(n926) );
  DFFR_X1 REG31_MY_CLK_r_REG157_S12 ( .D(REG31_n260), .CK(CLK), .RN(RST_n), 
        .Q(reg4[6]), .QN(n909) );
  DFFR_X1 REG31_MY_CLK_r_REG67_S14 ( .D(REG31_n262), .CK(CLK), .RN(RST_n), .Q(
        reg4[4]), .QN(n910) );
  DFFR_X1 REG31_MY_CLK_r_REG87_S17 ( .D(REG31_n264), .CK(CLK), .RN(RST_n), .Q(
        reg4[2]), .QN(n911) );
  DFFR_X1 REG31_MY_CLK_r_REG184_S6 ( .D(REG31_n254), .CK(CLK), .RN(RST_n), .Q(
        reg4[12]), .QN(n907) );
  DFFR_X1 REG31_MY_CLK_r_REG171_S10 ( .D(REG31_n256), .CK(CLK), .RN(RST_n), 
        .Q(reg4[10]), .QN(n912) );
  DFFR_X1 REG31_MY_CLK_r_REG141_S12 ( .D(REG31_n258), .CK(CLK), .RN(RST_n), 
        .Q(reg4[8]), .QN(n908) );
  DFFR_X1 REG41_MY_CLK_r_REG128_S15 ( .D(REG41_n263), .CK(CLK), .RN(RST_n), 
        .Q(reg5[3]), .QN(n933) );
  DFFR_X1 REG51_MY_CLK_r_REG69_S15 ( .D(REG51_n254), .CK(CLK), .RN(RST_n), 
        .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_) );
  DFFR_X1 REG51_MY_CLK_r_REG70_S15 ( .D(REG51_n255), .CK(CLK), .RN(RST_n), 
        .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_) );
  DFFR_X1 REG61_MY_CLK_r_REG192_S4 ( .D(REG61_n262), .CK(CLK), .RN(RST_n), .Q(
        reg7[5]), .QN(n897) );
  DFFR_X1 REG61_MY_CLK_r_REG187_S4 ( .D(REG61_n256), .CK(CLK), .RN(RST_n), .Q(
        reg7[11]), .QN(n913) );
  DFFR_X1 REG61_MY_CLK_r_REG18_S4 ( .D(REG61_n254), .CK(CLK), .RN(RST_n), .Q(
        reg7[13]), .QN(n914) );
  DFFR_X1 REG61_MY_CLK_r_REG34_S14 ( .D(REG61_n266), .CK(CLK), .RN(RST_n), .Q(
        reg7[1]), .QN(n900) );
  DFFR_X1 REG61_MY_CLK_r_REG31_S12 ( .D(REG61_n267), .CK(CLK), .RN(RST_n), .Q(
        reg7[0]), .QN(n882) );
  DFFR_X1 REG61_MY_CLK_r_REG174_S8 ( .D(REG61_n264), .CK(CLK), .RN(RST_n), .Q(
        reg7[3]), .QN(n896) );
  DFFR_X1 REG61_MY_CLK_r_REG189_S4 ( .D(REG61_n258), .CK(CLK), .RN(RST_n), .Q(
        reg7[9]), .QN(n899) );
  DFFR_X1 REG61_MY_CLK_r_REG191_S4 ( .D(REG61_n260), .CK(CLK), .RN(RST_n), .Q(
        reg7[7]), .QN(n898) );
  MUX2_X1 U235 ( .A(n70), .B(DIN[9]), .S(VIN), .Z(xin_in[9]) );
  MUX2_X1 U236 ( .A(n74), .B(DIN[8]), .S(VIN), .Z(xin_in[8]) );
  MUX2_X1 U237 ( .A(n75), .B(DIN[7]), .S(VIN), .Z(xin_in[7]) );
  MUX2_X1 U238 ( .A(n76), .B(DIN[6]), .S(VIN), .Z(xin_in[6]) );
  MUX2_X1 U239 ( .A(n77), .B(DIN[5]), .S(VIN), .Z(xin_in[5]) );
  MUX2_X1 U240 ( .A(n78), .B(DIN[4]), .S(VIN), .Z(xin_in[4]) );
  MUX2_X1 U241 ( .A(n79), .B(DIN[3]), .S(VIN), .Z(xin_in[3]) );
  MUX2_X1 U242 ( .A(n71), .B(DIN[2]), .S(VIN), .Z(xin_in[2]) );
  MUX2_X1 U243 ( .A(n72), .B(DIN[1]), .S(VIN), .Z(xin_in[1]) );
  MUX2_X1 U244 ( .A(n66), .B(DIN[13]), .S(VIN), .Z(xin_in[13]) );
  MUX2_X1 U245 ( .A(n67), .B(DIN[12]), .S(VIN), .Z(xin_in[12]) );
  MUX2_X1 U246 ( .A(n68), .B(DIN[11]), .S(VIN), .Z(xin_in[11]) );
  MUX2_X1 U247 ( .A(n69), .B(DIN[10]), .S(VIN), .Z(xin_in[10]) );
  MUX2_X1 U248 ( .A(n73), .B(DIN[0]), .S(VIN), .Z(xin_in[0]) );
  XOR2_X1 U249 ( .A(reg7[12]), .B(n279), .Z(SUB1_N12) );
  MUX2_X1 U250 ( .A(reg4_reg[0]), .B(reg5[0]), .S(VIN), .Z(REGISTER4_n266) );
  MUX2_X1 U251 ( .A(reg4_reg[1]), .B(reg5[1]), .S(VIN), .Z(REGISTER4_n265) );
  MUX2_X1 U252 ( .A(reg4_reg[2]), .B(reg5[2]), .S(VIN), .Z(REGISTER4_n264) );
  MUX2_X1 U254 ( .A(reg4_reg[4]), .B(reg5[4]), .S(VIN), .Z(REGISTER4_n262) );
  MUX2_X1 U256 ( .A(reg4_reg[6]), .B(reg5[6]), .S(VIN), .Z(REGISTER4_n260) );
  MUX2_X1 U258 ( .A(reg4_reg[8]), .B(reg5[8]), .S(VIN), .Z(REGISTER4_n258) );
  MUX2_X1 U260 ( .A(reg4_reg[10]), .B(reg5[10]), .S(VIN), .Z(REGISTER4_n256)
         );
  MUX2_X1 U262 ( .A(reg4_reg[12]), .B(reg5[12]), .S(VIN), .Z(REGISTER4_n254)
         );
  MUX2_X1 U264 ( .A(reg3_reg[0]), .B(reg3[0]), .S(VIN), .Z(REGISTER3_n266) );
  MUX2_X1 U266 ( .A(reg3_reg[2]), .B(reg3[2]), .S(VIN), .Z(REGISTER3_n264) );
  MUX2_X1 U268 ( .A(reg3_reg[4]), .B(reg3[4]), .S(VIN), .Z(REGISTER3_n262) );
  MUX2_X1 U269 ( .A(reg3_reg[5]), .B(reg3[5]), .S(VIN), .Z(REGISTER3_n261) );
  MUX2_X1 U270 ( .A(reg3_reg[6]), .B(reg3[6]), .S(VIN), .Z(REGISTER3_n260) );
  MUX2_X1 U271 ( .A(reg3_reg[7]), .B(reg3[7]), .S(VIN), .Z(REGISTER3_n259) );
  MUX2_X1 U272 ( .A(reg3_reg[8]), .B(reg3[8]), .S(VIN), .Z(REGISTER3_n258) );
  MUX2_X1 U273 ( .A(reg3_reg[9]), .B(reg3[9]), .S(VIN), .Z(REGISTER3_n257) );
  MUX2_X1 U274 ( .A(reg3_reg[10]), .B(reg3[10]), .S(VIN), .Z(REGISTER3_n256)
         );
  MUX2_X1 U275 ( .A(reg3_reg[11]), .B(reg3[11]), .S(VIN), .Z(REGISTER3_n255)
         );
  MUX2_X1 U276 ( .A(reg3_reg[12]), .B(reg3[12]), .S(VIN), .Z(REGISTER3_n254)
         );
  MUX2_X1 U277 ( .A(reg3_reg[13]), .B(reg3[13]), .S(VIN), .Z(REGISTER3_n253)
         );
  MUX2_X1 U278 ( .A(reg2_reg[0]), .B(reg2[0]), .S(VIN), .Z(REGISTER2_n266) );
  MUX2_X1 U279 ( .A(reg2_reg[1]), .B(reg2[1]), .S(VIN), .Z(REGISTER2_n265) );
  MUX2_X1 U280 ( .A(reg2_reg[2]), .B(reg2[2]), .S(VIN), .Z(REGISTER2_n264) );
  MUX2_X1 U281 ( .A(reg2_reg[4]), .B(reg2[4]), .S(VIN), .Z(REGISTER2_n262) );
  MUX2_X1 U282 ( .A(reg2_reg[5]), .B(reg2[5]), .S(VIN), .Z(REGISTER2_n261) );
  MUX2_X1 U283 ( .A(reg2_reg[6]), .B(reg2[6]), .S(VIN), .Z(REGISTER2_n260) );
  MUX2_X1 U284 ( .A(reg2_reg[7]), .B(reg2[7]), .S(VIN), .Z(REGISTER2_n259) );
  MUX2_X1 U285 ( .A(reg2_reg[8]), .B(reg2[8]), .S(VIN), .Z(REGISTER2_n258) );
  MUX2_X1 U286 ( .A(reg2_reg[9]), .B(reg2[9]), .S(VIN), .Z(REGISTER2_n257) );
  MUX2_X1 U287 ( .A(reg2_reg[10]), .B(reg2[10]), .S(VIN), .Z(REGISTER2_n256)
         );
  MUX2_X1 U288 ( .A(reg2_reg[11]), .B(reg2[11]), .S(VIN), .Z(REGISTER2_n255)
         );
  MUX2_X1 U289 ( .A(reg2_reg[12]), .B(reg2[12]), .S(VIN), .Z(REGISTER2_n254)
         );
  MUX2_X1 U290 ( .A(reg2_reg[13]), .B(reg2[13]), .S(VIN), .Z(REGISTER2_n253)
         );
  MUX2_X1 U291 ( .A(reg1_reg[3]), .B(w[3]), .S(VIN), .Z(REGISTER1_n263) );
  MUX2_X1 U292 ( .A(reg7[0]), .B(temp6[0]), .S(VIN), .Z(REG61_n267) );
  MUX2_X1 U293 ( .A(reg7[1]), .B(temp6[1]), .S(VIN), .Z(REG61_n266) );
  MUX2_X1 U294 ( .A(reg7[2]), .B(temp6[2]), .S(VIN), .Z(REG61_n265) );
  MUX2_X1 U295 ( .A(reg7[3]), .B(temp6[3]), .S(VIN), .Z(REG61_n264) );
  MUX2_X1 U296 ( .A(reg7[4]), .B(temp6[4]), .S(VIN), .Z(REG61_n263) );
  MUX2_X1 U297 ( .A(reg7[5]), .B(temp6[5]), .S(VIN), .Z(REG61_n262) );
  MUX2_X1 U298 ( .A(reg7[6]), .B(temp6[6]), .S(VIN), .Z(REG61_n261) );
  MUX2_X1 U299 ( .A(reg7[7]), .B(temp6[7]), .S(VIN), .Z(REG61_n260) );
  MUX2_X1 U300 ( .A(reg7[8]), .B(temp6[8]), .S(VIN), .Z(REG61_n259) );
  MUX2_X1 U301 ( .A(reg7[9]), .B(temp6[9]), .S(VIN), .Z(REG61_n258) );
  MUX2_X1 U302 ( .A(reg7[10]), .B(temp6[10]), .S(VIN), .Z(REG61_n257) );
  MUX2_X1 U303 ( .A(reg7[11]), .B(temp6[11]), .S(VIN), .Z(REG61_n256) );
  MUX2_X1 U304 ( .A(reg7[12]), .B(temp6[12]), .S(VIN), .Z(REG61_n255) );
  MUX2_X1 U306 ( .A(reg6[0]), .B(temp5[0]), .S(VIN), .Z(REG51_n266) );
  MUX2_X1 U307 ( .A(reg6[1]), .B(temp5[1]), .S(VIN), .Z(REG51_n265) );
  MUX2_X1 U308 ( .A(reg6[2]), .B(temp5[2]), .S(VIN), .Z(REG51_n264) );
  MUX2_X1 U309 ( .A(reg6[3]), .B(temp5[3]), .S(VIN), .Z(REG51_n263) );
  MUX2_X1 U310 ( .A(reg6[4]), .B(temp5[4]), .S(VIN), .Z(REG51_n262) );
  MUX2_X1 U311 ( .A(reg6[5]), .B(temp5[5]), .S(VIN), .Z(REG51_n261) );
  MUX2_X1 U312 ( .A(reg6[6]), .B(temp5[6]), .S(VIN), .Z(REG51_n260) );
  MUX2_X1 U313 ( .A(reg6[7]), .B(temp5[7]), .S(VIN), .Z(REG51_n259) );
  MUX2_X1 U314 ( .A(reg6[8]), .B(temp5[8]), .S(VIN), .Z(REG51_n258) );
  MUX2_X1 U315 ( .A(reg6[9]), .B(temp5[9]), .S(VIN), .Z(REG51_n257) );
  MUX2_X1 U316 ( .A(reg6[10]), .B(temp5[10]), .S(VIN), .Z(REG51_n256) );
  MUX2_X1 U320 ( .A(mul4_reg[0]), .B(temp4[0]), .S(VIN), .Z(REG4_1_n266) );
  MUX2_X1 U321 ( .A(mul4_reg[1]), .B(temp4[1]), .S(VIN), .Z(REG4_1_n265) );
  MUX2_X1 U322 ( .A(mul4_reg[2]), .B(temp4[2]), .S(VIN), .Z(REG4_1_n264) );
  MUX2_X1 U323 ( .A(mul4_reg[3]), .B(temp4[3]), .S(VIN), .Z(REG4_1_n263) );
  MUX2_X1 U324 ( .A(mul4_reg[4]), .B(temp4[4]), .S(VIN), .Z(REG4_1_n262) );
  MUX2_X1 U325 ( .A(mul4_reg[5]), .B(temp4[5]), .S(VIN), .Z(REG4_1_n261) );
  MUX2_X1 U326 ( .A(mul4_reg[6]), .B(temp4[6]), .S(VIN), .Z(REG4_1_n260) );
  MUX2_X1 U327 ( .A(mul4_reg[7]), .B(temp4[7]), .S(VIN), .Z(REG4_1_n259) );
  MUX2_X1 U328 ( .A(mul4_reg[8]), .B(temp4[8]), .S(VIN), .Z(REG4_1_n258) );
  MUX2_X1 U329 ( .A(mul4_reg[9]), .B(temp4[9]), .S(VIN), .Z(REG4_1_n257) );
  MUX2_X1 U330 ( .A(mul4_reg[10]), .B(temp4[10]), .S(VIN), .Z(REG4_1_n256) );
  MUX2_X1 U331 ( .A(mul4_reg[11]), .B(temp4[11]), .S(VIN), .Z(REG4_1_n255) );
  MUX2_X1 U334 ( .A(mul3_reg[0]), .B(temp3[0]), .S(VIN), .Z(REG3_1_n267) );
  MUX2_X1 U335 ( .A(mul3_reg[1]), .B(temp3[1]), .S(VIN), .Z(REG3_1_n266) );
  MUX2_X1 U336 ( .A(mul3_reg[2]), .B(temp3[2]), .S(VIN), .Z(REG3_1_n265) );
  MUX2_X1 U337 ( .A(mul3_reg[3]), .B(temp3[3]), .S(VIN), .Z(REG3_1_n264) );
  MUX2_X1 U338 ( .A(mul3_reg[4]), .B(temp3[4]), .S(VIN), .Z(REG3_1_n263) );
  MUX2_X1 U339 ( .A(mul3_reg[5]), .B(temp3[5]), .S(VIN), .Z(REG3_1_n262) );
  MUX2_X1 U340 ( .A(mul3_reg[6]), .B(temp3[6]), .S(VIN), .Z(REG3_1_n261) );
  MUX2_X1 U341 ( .A(mul3_reg[7]), .B(temp3[7]), .S(VIN), .Z(REG3_1_n260) );
  MUX2_X1 U342 ( .A(mul3_reg[8]), .B(temp3[8]), .S(VIN), .Z(REG3_1_n259) );
  MUX2_X1 U343 ( .A(mul3_reg[9]), .B(temp3[9]), .S(VIN), .Z(REG3_1_n258) );
  MUX2_X1 U344 ( .A(mul3_reg[10]), .B(temp3[10]), .S(VIN), .Z(REG3_1_n257) );
  MUX2_X1 U345 ( .A(mul3_reg[11]), .B(temp3[11]), .S(VIN), .Z(REG3_1_n256) );
  MUX2_X1 U346 ( .A(mul3_reg[12]), .B(temp3[12]), .S(VIN), .Z(REG3_1_n255) );
  MUX2_X1 U348 ( .A(mul2_reg[0]), .B(temp2[0]), .S(VIN), .Z(REG2_1_n270) );
  MUX2_X1 U349 ( .A(mul2_reg[1]), .B(temp2[1]), .S(VIN), .Z(REG2_1_n269) );
  MUX2_X1 U350 ( .A(mul2_reg[2]), .B(temp2[2]), .S(VIN), .Z(REG2_1_n268) );
  MUX2_X1 U351 ( .A(mul2_reg[3]), .B(temp2[3]), .S(VIN), .Z(REG2_1_n267) );
  MUX2_X1 U352 ( .A(mul2_reg[4]), .B(temp2[4]), .S(VIN), .Z(REG2_1_n266) );
  MUX2_X1 U353 ( .A(mul2_reg[5]), .B(temp2[5]), .S(VIN), .Z(REG2_1_n265) );
  MUX2_X1 U354 ( .A(mul2_reg[6]), .B(temp2[6]), .S(VIN), .Z(REG2_1_n264) );
  MUX2_X1 U355 ( .A(mul2_reg[7]), .B(temp2[7]), .S(VIN), .Z(REG2_1_n263) );
  MUX2_X1 U356 ( .A(mul2_reg[8]), .B(temp2[8]), .S(VIN), .Z(REG2_1_n262) );
  MUX2_X1 U357 ( .A(mul2_reg[9]), .B(temp2[9]), .S(VIN), .Z(REG2_1_n261) );
  MUX2_X1 U358 ( .A(mul2_reg[10]), .B(temp2[10]), .S(VIN), .Z(REG2_1_n260) );
  MUX2_X1 U360 ( .A(mul2_reg[12]), .B(temp2[12]), .S(VIN), .Z(REG2_1_n258) );
  MUX2_X1 U361 ( .A(mul1_reg[0]), .B(temp1[0]), .S(VIN), .Z(REG1_1_n267) );
  MUX2_X1 U362 ( .A(mul1_reg[1]), .B(temp1[1]), .S(VIN), .Z(REG1_1_n266) );
  MUX2_X1 U363 ( .A(mul1_reg[2]), .B(temp1[2]), .S(VIN), .Z(REG1_1_n265) );
  MUX2_X1 U364 ( .A(mul1_reg[3]), .B(temp1[3]), .S(VIN), .Z(REG1_1_n264) );
  MUX2_X1 U365 ( .A(mul1_reg[4]), .B(temp1[4]), .S(VIN), .Z(REG1_1_n263) );
  MUX2_X1 U366 ( .A(mul1_reg[5]), .B(temp1[5]), .S(VIN), .Z(REG1_1_n262) );
  MUX2_X1 U367 ( .A(mul1_reg[6]), .B(temp1[6]), .S(VIN), .Z(REG1_1_n261) );
  MUX2_X1 U368 ( .A(mul1_reg[7]), .B(temp1[7]), .S(VIN), .Z(REG1_1_n260) );
  MUX2_X1 U369 ( .A(mul1_reg[8]), .B(temp1[8]), .S(VIN), .Z(REG1_1_n259) );
  MUX2_X1 U370 ( .A(mul1_reg[9]), .B(temp1[9]), .S(VIN), .Z(REG1_1_n258) );
  MUX2_X1 U371 ( .A(mul1_reg[10]), .B(temp1[10]), .S(VIN), .Z(REG1_1_n257) );
  MUX2_X1 U372 ( .A(mul1_reg[11]), .B(temp1[11]), .S(VIN), .Z(REG1_1_n256) );
  MUX2_X1 U373 ( .A(mul1_reg[12]), .B(temp1[12]), .S(VIN), .Z(REG1_1_n255) );
  DFFR_X1 REG31_MY_CLK_r_REG117_S17 ( .D(REG31_n266), .CK(CLK), .RN(RST_n), 
        .Q(reg4[0]), .QN(n906) );
  DFFR_X1 REG31_MY_CLK_r_REG196_S4 ( .D(REG31_n253), .CK(CLK), .RN(RST_n), .Q(
        reg4[13]), .QN(n903) );
  DFFR_X1 REG31_MY_CLK_r_REG149_S12 ( .D(REG31_n259), .CK(CLK), .RN(RST_n), 
        .Q(reg4[7]), .QN(n904) );
  DFFR_X1 REG31_MY_CLK_r_REG178_S8 ( .D(REG31_n255), .CK(CLK), .RN(RST_n), .Q(
        reg4[11]), .QN(n902) );
  DFFR_X1 REG31_MY_CLK_r_REG133_S12 ( .D(REG31_n257), .CK(CLK), .RN(RST_n), 
        .Q(reg4[9]), .QN(n901) );
  DFFR_X1 REG11_MY_CLK_r_REG17_S3 ( .D(REG11_n254), .CK(CLK), .RN(RST_n), .Q(
        reg2[13]), .QN(n887) );
  DFFR_X1 REG11_MY_CLK_r_REG161_S11 ( .D(REG11_n262), .CK(CLK), .RN(RST_n), 
        .Q(reg2[5]), .QN(n886) );
  DFFR_X1 REG11_MY_CLK_r_REG145_S11 ( .D(REG11_n260), .CK(CLK), .RN(RST_n), 
        .Q(reg2[7]), .QN(n885) );
  DFFR_X1 REG11_MY_CLK_r_REG30_S11 ( .D(REG11_n258), .CK(CLK), .RN(RST_n), .Q(
        reg2[9]), .QN(n884) );
  DFFR_X1 REG11_MY_CLK_r_REG24_S7 ( .D(REG11_n256), .CK(CLK), .RN(RST_n), .Q(
        reg2[11]), .QN(n883) );
  NAND2_X1 U69 ( .A1(n268), .A2(n897), .ZN(n267) );
  NAND2_X1 U66 ( .A1(n263), .A2(n898), .ZN(n262) );
  NAND2_X1 U63 ( .A1(n260), .A2(n899), .ZN(n282) );
  NOR2_X1 U60 ( .A1(reg7[10]), .A2(n282), .ZN(n280) );
  NAND2_X1 U57 ( .A1(n280), .A2(n913), .ZN(n279) );
  NOR2_X1 U56 ( .A1(n279), .A2(reg7[12]), .ZN(n278) );
  XNOR2_X1 U55 ( .A(n278), .B(reg7[13]), .ZN(SUB1_N13) );
  XNOR2_X1 U59 ( .A(reg7[11]), .B(n280), .ZN(SUB1_N11) );
  NOR2_X1 U62 ( .A1(reg7[10]), .A2(reg7[9]), .ZN(n283) );
  AOI22_X1 U61 ( .A1(n282), .A2(reg7[10]), .B1(n260), .B2(n283), .ZN(SUB1_N10)
         );
  AOI22_X1 U39 ( .A1(reg7[9]), .A2(n259), .B1(n260), .B2(n899), .ZN(SUB1_N9)
         );
  NOR2_X1 U42 ( .A1(reg7[8]), .A2(reg7[7]), .ZN(n264) );
  AOI22_X1 U41 ( .A1(n262), .A2(reg7[8]), .B1(n263), .B2(n264), .ZN(SUB1_N8)
         );
  AOI22_X1 U43 ( .A1(n263), .A2(n898), .B1(reg7[7]), .B2(n266), .ZN(SUB1_N7)
         );
  NOR2_X1 U46 ( .A1(reg7[6]), .A2(reg7[5]), .ZN(n269) );
  AOI22_X1 U45 ( .A1(n267), .A2(reg7[6]), .B1(n268), .B2(n269), .ZN(SUB1_N6)
         );
  AOI22_X1 U47 ( .A1(n268), .A2(n897), .B1(reg7[5]), .B2(n271), .ZN(SUB1_N5)
         );
  NOR2_X1 U50 ( .A1(reg7[4]), .A2(reg7[3]), .ZN(n274) );
  AOI22_X1 U49 ( .A1(n272), .A2(reg7[4]), .B1(n273), .B2(n274), .ZN(SUB1_N4)
         );
  AOI22_X1 U51 ( .A1(n273), .A2(n896), .B1(reg7[3]), .B2(n276), .ZN(SUB1_N3)
         );
  NOR2_X1 U54 ( .A1(reg7[1]), .A2(reg7[0]), .ZN(n277) );
  XNOR2_X1 U53 ( .A(n277), .B(reg7[2]), .ZN(SUB1_N2) );
  AOI22_X1 U75 ( .A1(reg7[0]), .A2(reg7[1]), .B1(n900), .B2(n882), .ZN(SUB1_N1) );
  NAND2_X1 U233 ( .A1(VIN), .A2(w[13]), .ZN(n312) );
  OAI21_X1 U232 ( .B1(VIN), .B2(n887), .A(n312), .ZN(REG11_n254) );
  NAND2_X1 U105 ( .A1(reg1_reg[13]), .A2(n942), .ZN(n313) );
  NAND2_X1 U104 ( .A1(n312), .A2(n313), .ZN(REGISTER1_n253) );
  NAND2_X1 U230 ( .A1(VIN), .A2(w[12]), .ZN(n310) );
  OAI21_X1 U229 ( .B1(VIN), .B2(n890), .A(n310), .ZN(REG11_n255) );
  NAND2_X1 U103 ( .A1(reg1_reg[12]), .A2(n940), .ZN(n311) );
  NAND2_X1 U102 ( .A1(n310), .A2(n311), .ZN(REGISTER1_n254) );
  NAND2_X1 U227 ( .A1(VIN), .A2(w[11]), .ZN(n308) );
  OAI21_X1 U226 ( .B1(VIN), .B2(n883), .A(n308), .ZN(REG11_n256) );
  NAND2_X1 U101 ( .A1(reg1_reg[11]), .A2(n940), .ZN(n309) );
  NAND2_X1 U100 ( .A1(n308), .A2(n309), .ZN(REGISTER1_n255) );
  NAND2_X1 U224 ( .A1(VIN), .A2(w[10]), .ZN(n306) );
  OAI21_X1 U223 ( .B1(VIN), .B2(n891), .A(n306), .ZN(REG11_n257) );
  NAND2_X1 U99 ( .A1(reg1_reg[10]), .A2(n942), .ZN(n307) );
  NAND2_X1 U98 ( .A1(n306), .A2(n307), .ZN(REGISTER1_n256) );
  NAND2_X1 U221 ( .A1(VIN), .A2(w[9]), .ZN(n304) );
  OAI21_X1 U220 ( .B1(VIN), .B2(n884), .A(n304), .ZN(REG11_n258) );
  NAND2_X1 U97 ( .A1(reg1_reg[9]), .A2(n942), .ZN(n305) );
  NAND2_X1 U96 ( .A1(n304), .A2(n305), .ZN(REGISTER1_n257) );
  NAND2_X1 U218 ( .A1(VIN), .A2(w[8]), .ZN(n302) );
  OAI21_X1 U217 ( .B1(VIN), .B2(n892), .A(n302), .ZN(REG11_n259) );
  NAND2_X1 U95 ( .A1(reg1_reg[8]), .A2(n942), .ZN(n303) );
  NAND2_X1 U94 ( .A1(n302), .A2(n303), .ZN(REGISTER1_n258) );
  NAND2_X1 U215 ( .A1(VIN), .A2(w[7]), .ZN(n300) );
  OAI21_X1 U214 ( .B1(VIN), .B2(n885), .A(n300), .ZN(REG11_n260) );
  NAND2_X1 U93 ( .A1(reg1_reg[7]), .A2(n940), .ZN(n301) );
  NAND2_X1 U92 ( .A1(n300), .A2(n301), .ZN(REGISTER1_n259) );
  NAND2_X1 U212 ( .A1(VIN), .A2(w[6]), .ZN(n298) );
  OAI21_X1 U211 ( .B1(VIN), .B2(n893), .A(n298), .ZN(REG11_n261) );
  NAND2_X1 U91 ( .A1(reg1_reg[6]), .A2(n941), .ZN(n299) );
  NAND2_X1 U90 ( .A1(n298), .A2(n299), .ZN(REGISTER1_n260) );
  NAND2_X1 U209 ( .A1(VIN), .A2(w[5]), .ZN(n296) );
  OAI21_X1 U208 ( .B1(VIN), .B2(n886), .A(n296), .ZN(REG11_n262) );
  NAND2_X1 U89 ( .A1(reg1_reg[5]), .A2(n942), .ZN(n297) );
  NAND2_X1 U88 ( .A1(n296), .A2(n297), .ZN(REGISTER1_n261) );
  NAND2_X1 U206 ( .A1(VIN), .A2(w[4]), .ZN(n294) );
  OAI21_X1 U205 ( .B1(VIN), .B2(n894), .A(n294), .ZN(REG11_n263) );
  NAND2_X1 U87 ( .A1(reg1_reg[4]), .A2(n940), .ZN(n295) );
  NAND2_X1 U86 ( .A1(n294), .A2(n295), .ZN(REGISTER1_n262) );
  OAI22_X1 U125 ( .A1(n941), .A2(reg4[9]), .B1(reg5[9]), .B2(VIN), .ZN(n324)
         );
  OAI22_X1 U129 ( .A1(n941), .A2(reg4[11]), .B1(reg5[11]), .B2(VIN), .ZN(n326)
         );
  OAI22_X1 U121 ( .A1(n941), .A2(reg4[7]), .B1(reg5[7]), .B2(VIN), .ZN(n322)
         );
  OAI22_X1 U133 ( .A1(n941), .A2(reg4[13]), .B1(reg5[13]), .B2(VIN), .ZN(n328)
         );
  OAI22_X1 U119 ( .A1(n941), .A2(reg4[6]), .B1(reg5[6]), .B2(VIN), .ZN(n321)
         );
  OAI22_X1 U123 ( .A1(n941), .A2(reg4[8]), .B1(reg5[8]), .B2(VIN), .ZN(n323)
         );
  OAI22_X1 U127 ( .A1(n941), .A2(reg4[10]), .B1(reg5[10]), .B2(VIN), .ZN(n325)
         );
  OAI22_X1 U131 ( .A1(n941), .A2(reg4[12]), .B1(reg5[12]), .B2(VIN), .ZN(n327)
         );
  OAI22_X1 U111 ( .A1(n941), .A2(reg4[2]), .B1(reg5[2]), .B2(VIN), .ZN(n316)
         );
  OAI22_X1 U115 ( .A1(n941), .A2(reg4[4]), .B1(reg5[4]), .B2(VIN), .ZN(n319)
         );
  OAI22_X1 U107 ( .A1(n941), .A2(reg4[0]), .B1(reg5[0]), .B2(VIN), .ZN(n314)
         );
  OAI22_X1 U117 ( .A1(n941), .A2(reg4[5]), .B1(reg5[5]), .B2(VIN), .ZN(n320)
         );
  AOI22_X1 U194 ( .A1(VIN), .A2(w[3]), .B1(reg2[3]), .B2(n941), .ZN(REG11_n64)
         );
  NAND2_X1 U200 ( .A1(VIN), .A2(w[1]), .ZN(n290) );
  NAND2_X1 U83 ( .A1(reg1_reg[1]), .A2(n941), .ZN(n291) );
  NAND2_X1 U82 ( .A1(n290), .A2(n291), .ZN(REGISTER1_n265) );
  NAND2_X1 U203 ( .A1(VIN), .A2(w[2]), .ZN(n292) );
  OAI21_X1 U202 ( .B1(VIN), .B2(n895), .A(n292), .ZN(REG11_n264) );
  NAND2_X1 U85 ( .A1(reg1_reg[2]), .A2(n942), .ZN(n293) );
  NAND2_X1 U84 ( .A1(n292), .A2(n293), .ZN(REGISTER1_n264) );
  NAND2_X1 U81 ( .A1(reg1_reg[0]), .A2(n940), .ZN(n289) );
  NAND2_X1 U80 ( .A1(n288), .A2(n289), .ZN(REGISTER1_n266) );
  NAND2_X1 U79 ( .A1(reg2_reg[3]), .A2(n940), .ZN(n287) );
  OAI21_X1 U171 ( .B1(VIN), .B2(n919), .A(n286), .ZN(REG21_n263) );
  OAI21_X1 U199 ( .B1(VIN), .B2(n888), .A(n290), .ZN(REG11_n265) );
  OAI21_X1 U196 ( .B1(VIN), .B2(p11_mult_21_n693), .A(n288), .ZN(REG11_n266)
         );
  AOI22_X1 U186 ( .A1(VIN), .A2(n891), .B1(n923), .B2(n941), .ZN(REG21_n256)
         );
  AOI22_X1 U180 ( .A1(VIN), .A2(n885), .B1(n926), .B2(n941), .ZN(REG21_n259)
         );
  AOI22_X1 U182 ( .A1(VIN), .A2(n892), .B1(n925), .B2(n940), .ZN(REG21_n258)
         );
  AOI22_X1 U188 ( .A1(VIN), .A2(n883), .B1(n922), .B2(n942), .ZN(REG21_n255)
         );
  AOI22_X1 U165 ( .A1(VIN), .A2(p11_mult_21_n693), .B1(n932), .B2(n940), .ZN(
        REG21_n266) );
  AOI22_X1 U169 ( .A1(VIN), .A2(n895), .B1(n930), .B2(n940), .ZN(REG21_n264)
         );
  AOI22_X1 U160 ( .A1(VIN), .A2(n887), .B1(n903), .B2(n942), .ZN(REG31_n253)
         );
  AOI22_X1 U150 ( .A1(VIN), .A2(n892), .B1(n908), .B2(n942), .ZN(REG31_n258)
         );
  AOI22_X1 U154 ( .A1(VIN), .A2(n891), .B1(n912), .B2(n940), .ZN(REG31_n256)
         );
  AOI22_X1 U192 ( .A1(VIN), .A2(n887), .B1(n920), .B2(n940), .ZN(REG21_n253)
         );
  AOI22_X1 U176 ( .A1(VIN), .A2(n886), .B1(n928), .B2(n940), .ZN(REG21_n261)
         );
  AOI22_X1 U142 ( .A1(VIN), .A2(n894), .B1(n910), .B2(n942), .ZN(REG31_n262)
         );
  AOI22_X1 U146 ( .A1(VIN), .A2(n893), .B1(n909), .B2(n942), .ZN(REG31_n260)
         );
  AOI22_X1 U144 ( .A1(VIN), .A2(n886), .B1(p10_mult_21_n1046), .B2(n942), .ZN(
        REG31_n261) );
  AOI22_X1 U134 ( .A1(VIN), .A2(p11_mult_21_n693), .B1(n906), .B2(n940), .ZN(
        REG31_n266) );
  AOI22_X1 U184 ( .A1(VIN), .A2(n884), .B1(n924), .B2(n941), .ZN(REG21_n257)
         );
  AOI22_X1 U178 ( .A1(VIN), .A2(n893), .B1(n927), .B2(n941), .ZN(REG21_n260)
         );
  AOI22_X1 U156 ( .A1(VIN), .A2(n883), .B1(n902), .B2(n942), .ZN(REG31_n255)
         );
  AOI22_X1 U136 ( .A1(VIN), .A2(n888), .B1(n905), .B2(n942), .ZN(REG31_n265)
         );
  AOI22_X1 U174 ( .A1(VIN), .A2(n894), .B1(n929), .B2(n940), .ZN(REG21_n262)
         );
  AOI22_X1 U190 ( .A1(VIN), .A2(n890), .B1(n921), .B2(n940), .ZN(REG21_n254)
         );
  AOI22_X1 U167 ( .A1(VIN), .A2(n888), .B1(n931), .B2(n940), .ZN(REG21_n265)
         );
  AOI22_X1 U148 ( .A1(VIN), .A2(n885), .B1(n904), .B2(n942), .ZN(REG31_n259)
         );
  AOI22_X1 U152 ( .A1(VIN), .A2(n884), .B1(n901), .B2(n940), .ZN(REG31_n257)
         );
  AOI22_X1 U138 ( .A1(VIN), .A2(n895), .B1(n911), .B2(n940), .ZN(REG31_n264)
         );
  AOI22_X1 U158 ( .A1(VIN), .A2(n890), .B1(n907), .B2(n940), .ZN(REG31_n254)
         );
  AOI22_X1 U112 ( .A1(VIN), .A2(n889), .B1(n933), .B2(n940), .ZN(REG41_n263)
         );
  NAND2_X1 U38 ( .A1(n30), .A2(n942), .ZN(n185) );
  NAND2_X1 U163 ( .A1(n940), .A2(mul2_reg[13]), .ZN(REG2_1_n272) );
  NAND2_X1 U172 ( .A1(VIN), .A2(reg2[3]), .ZN(n286) );
  MUX2_X1 U265 ( .A(reg3_reg[1]), .B(reg3[1]), .S(VIN), .Z(REGISTER3_n265) );
  MUX2_X1 U259 ( .A(reg4_reg[9]), .B(reg5[9]), .S(VIN), .Z(REGISTER4_n257) );
  MUX2_X1 U257 ( .A(reg4_reg[7]), .B(reg5[7]), .S(VIN), .Z(REGISTER4_n259) );
  MUX2_X1 U261 ( .A(reg4_reg[11]), .B(reg5[11]), .S(VIN), .Z(REGISTER4_n255)
         );
  MUX2_X1 U263 ( .A(reg4_reg[13]), .B(reg5[13]), .S(VIN), .Z(REGISTER4_n253)
         );
  MUX2_X1 U267 ( .A(reg3_reg[3]), .B(reg3[3]), .S(VIN), .Z(REGISTER3_n263) );
  MUX2_X1 U255 ( .A(reg4_reg[5]), .B(reg5[5]), .S(VIN), .Z(REGISTER4_n261) );
  MUX2_X1 U253 ( .A(reg4_reg[3]), .B(reg5[3]), .S(VIN), .Z(REGISTER4_n263) );
  NAND2_X1 U72 ( .A1(n273), .A2(n896), .ZN(n272) );
  NOR3_X1 U74 ( .A1(reg7[0]), .A2(reg7[2]), .A3(reg7[1]), .ZN(n273) );
  NOR2_X1 U68 ( .A1(reg7[6]), .A2(n267), .ZN(n263) );
  NOR2_X1 U65 ( .A1(reg7[8]), .A2(n262), .ZN(n260) );
  NOR2_X1 U71 ( .A1(reg7[4]), .A2(n272), .ZN(n268) );
  INV_X1 U40 ( .A(n260), .ZN(n259) );
  INV_X1 U44 ( .A(n263), .ZN(n266) );
  INV_X1 U48 ( .A(n268), .ZN(n271) );
  INV_X1 U52 ( .A(n273), .ZN(n276) );
  OR2_X1 U164 ( .A1(REG2_1_n271), .A2(REG2_1_n92), .ZN(mul2_reg[13]) );
  INV_X1 U124 ( .A(n324), .ZN(REG41_n257) );
  INV_X1 U128 ( .A(n326), .ZN(REG41_n255) );
  INV_X1 U120 ( .A(n322), .ZN(REG41_n259) );
  INV_X1 U132 ( .A(n328), .ZN(REG41_n253) );
  INV_X1 U118 ( .A(n321), .ZN(REG41_n260) );
  INV_X1 U122 ( .A(n323), .ZN(REG41_n258) );
  INV_X1 U126 ( .A(n325), .ZN(REG41_n256) );
  INV_X1 U130 ( .A(n327), .ZN(REG41_n254) );
  INV_X1 U110 ( .A(n316), .ZN(REG41_n264) );
  INV_X1 U114 ( .A(n319), .ZN(REG41_n262) );
  INV_X1 U106 ( .A(n314), .ZN(REG41_n266) );
  INV_X1 U116 ( .A(n320), .ZN(REG41_n261) );
  INV_X1 U108 ( .A(n315), .ZN(REG41_n265) );
  INV_X1 p6_mult_21_U717 ( .A(p6_mult_21_n267), .ZN(p6_mult_21_n827) );
  INV_X1 p6_mult_21_U718 ( .A(p6_mult_21_n258), .ZN(p6_mult_21_n826) );
  AND3_X1 p6_mult_21_U413 ( .A1(p6_mult_21_n678), .A2(p6_mult_21_n679), .A3(
        p6_mult_21_n680), .ZN(p6_mult_21_n825) );
  INV_X1 p6_mult_21_U720 ( .A(p6_mult_21_n285), .ZN(p6_mult_21_n831) );
  INV_X1 p6_mult_21_U721 ( .A(p6_mult_21_n278), .ZN(p6_mult_21_n830) );
  AND3_X1 p6_mult_21_U410 ( .A1(p6_mult_21_n659), .A2(p6_mult_21_n660), .A3(
        p6_mult_21_n661), .ZN(p6_mult_21_n829) );
  INV_X1 p6_mult_21_U735 ( .A(p6_mult_21_n842), .ZN(p6_mult_21_n844) );
  INV_X1 p6_mult_21_U729 ( .A(B0[0]), .ZN(p6_mult_21_n722) );
  OR2_X1 p6_mult_21_U670 ( .A1(p6_mult_21_n817), .A2(p6_mult_21_n818), .ZN(
        p6_mult_21_n243) );
  INV_X1 p6_mult_21_U502 ( .A(p6_mult_21_n703), .ZN(p6_mult_21_n408) );
  INV_X1 p6_mult_21_U529 ( .A(p6_mult_21_n720), .ZN(p6_mult_21_n394) );
  INV_X1 p6_mult_21_U677 ( .A(p6_mult_21_n231), .ZN(p6_mult_21_n232) );
  INV_X1 p6_mult_21_U424 ( .A(p6_mult_21_n837), .ZN(p6_mult_21_n707) );
  INV_X1 p6_mult_21_U681 ( .A(p6_mult_21_n209), .ZN(p6_mult_21_n210) );
  INV_X1 p6_mult_21_U553 ( .A(p6_mult_21_n738), .ZN(p6_mult_21_n380) );
  NAND2_X1 p6_mult_21_U453 ( .A1(p6_mult_21_n723), .A2(p6_mult_21_n819), .ZN(
        p6_mult_21_n725) );
  INV_X1 p6_mult_21_U686 ( .A(p6_mult_21_n191), .ZN(p6_mult_21_n192) );
  INV_X1 p6_mult_21_U580 ( .A(p6_mult_21_n755), .ZN(p6_mult_21_n366) );
  NAND2_X1 p6_mult_21_U689 ( .A1(p6_mult_21_n740), .A2(p6_mult_21_n821), .ZN(
        p6_mult_21_n742) );
  INV_X1 p6_mult_21_U693 ( .A(p6_mult_21_n177), .ZN(p6_mult_21_n178) );
  INV_X1 p6_mult_21_U607 ( .A(p6_mult_21_n772), .ZN(p6_mult_21_n352) );
  NAND2_X1 p6_mult_21_U696 ( .A1(p6_mult_21_n757), .A2(p6_mult_21_n822), .ZN(
        p6_mult_21_n759) );
  INV_X1 p6_mult_21_U700 ( .A(p6_mult_21_n167), .ZN(p6_mult_21_n168) );
  INV_X1 p6_mult_21_U709 ( .A(p6_mult_21_n791), .ZN(p6_mult_21_n687) );
  INV_X1 p6_mult_21_U710 ( .A(p6_mult_21_n793), .ZN(p6_mult_21_n686) );
  INV_X1 p6_mult_21_U631 ( .A(p6_mult_21_n789), .ZN(p6_mult_21_n338) );
  INV_X1 p6_mult_21_U657 ( .A(p6_mult_21_n806), .ZN(p6_mult_21_n805) );
  NAND2_X1 p6_mult_21_U703 ( .A1(p6_mult_21_n774), .A2(p6_mult_21_n823), .ZN(
        p6_mult_21_n776) );
  NAND2_X1 p6_mult_21_U724 ( .A1(p6_mult_21_n707), .A2(p6_mult_21_n838), .ZN(
        p6_mult_21_n706) );
  NAND2_X1 p6_mult_21_U711 ( .A1(p6_mult_21_n791), .A2(p6_mult_21_n824), .ZN(
        p6_mult_21_n793) );
  NAND2_X1 p6_mult_21_U464 ( .A1(p6_mult_21_n246), .A2(p6_mult_21_n257), .ZN(
        p6_mult_21_n674) );
  NAND2_X1 p6_mult_21_U463 ( .A1(p6_mult_21_n149), .A2(p6_mult_21_n257), .ZN(
        p6_mult_21_n673) );
  OAI222_X1 p6_mult_21_U716 ( .A1(p6_mult_21_n825), .A2(p6_mult_21_n826), .B1(
        p6_mult_21_n825), .B2(p6_mult_21_n827), .C1(p6_mult_21_n827), .C2(
        p6_mult_21_n826), .ZN(p6_mult_21_n149) );
  NAND2_X1 p6_mult_21_U471 ( .A1(p6_mult_21_n277), .A2(p6_mult_21_n268), .ZN(
        p6_mult_21_n680) );
  OAI22_X1 p6_mult_21_U521 ( .A1(p6_mult_21_n715), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n716), .ZN(p6_mult_21_n398) );
  OAI22_X1 p6_mult_21_U564 ( .A1(p6_mult_21_n746), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n747), .ZN(p6_mult_21_n374) );
  OAI222_X1 p6_mult_21_U719 ( .A1(p6_mult_21_n829), .A2(p6_mult_21_n830), .B1(
        p6_mult_21_n829), .B2(p6_mult_21_n831), .C1(p6_mult_21_n831), .C2(
        p6_mult_21_n830), .ZN(p6_mult_21_n828) );
  OAI22_X1 p6_mult_21_U494 ( .A1(p6_mult_21_n698), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n699), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n412) );
  NOR2_X1 p6_mult_21_U609 ( .A1(p6_mult_21_n722), .A2(p6_mult_21_n774), .ZN(
        p6_mult_21_n351) );
  OAI22_X1 p6_mult_21_U562 ( .A1(p6_mult_21_n745), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n746), .ZN(p6_mult_21_n375) );
  XNOR2_X1 p6_mult_21_U565 ( .A(B0[4]), .B(reg1_reg[7]), .ZN(p6_mult_21_n746)
         );
  OAI22_X1 p6_mult_21_U519 ( .A1(p6_mult_21_n714), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n715), .ZN(p6_mult_21_n399) );
  OAI22_X1 p6_mult_21_U585 ( .A1(p6_mult_21_n760), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n761), .ZN(p6_mult_21_n363) );
  NAND2_X1 p6_mult_21_U446 ( .A1(p6_mult_21_n293), .A2(p6_mult_21_n286), .ZN(
        p6_mult_21_n661) );
  NAND2_X1 p6_mult_21_U445 ( .A1(p6_mult_21_n635), .A2(p6_mult_21_n293), .ZN(
        p6_mult_21_n660) );
  NAND2_X1 p6_mult_21_U444 ( .A1(p6_mult_21_n635), .A2(p6_mult_21_n286), .ZN(
        p6_mult_21_n659) );
  OAI22_X1 p6_mult_21_U492 ( .A1(p6_mult_21_n697), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n698), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n413) );
  XNOR2_X1 p6_mult_21_U495 ( .A(B0[9]), .B(reg1_reg[1]), .ZN(p6_mult_21_n698)
         );
  XNOR2_X1 p6_mult_21_U586 ( .A(B0[1]), .B(reg1_reg[9]), .ZN(p6_mult_21_n760)
         );
  OAI22_X1 p6_mult_21_U517 ( .A1(p6_mult_21_n713), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n714), .ZN(p6_mult_21_n400) );
  XNOR2_X1 p6_mult_21_U543 ( .A(B0[5]), .B(reg1_reg[5]), .ZN(p6_mult_21_n730)
         );
  OAI22_X1 p6_mult_21_U560 ( .A1(p6_mult_21_n744), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n745), .ZN(p6_mult_21_n376) );
  XNOR2_X1 p6_mult_21_U563 ( .A(B0[3]), .B(reg1_reg[7]), .ZN(p6_mult_21_n745)
         );
  NAND2_X1 p6_mult_21_U419 ( .A1(p6_mult_21_n299), .A2(p6_mult_21_n294), .ZN(
        p6_mult_21_n643) );
  OAI22_X1 p6_mult_21_U515 ( .A1(p6_mult_21_n712), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n713), .ZN(p6_mult_21_n401) );
  OAI22_X1 p6_mult_21_U558 ( .A1(p6_mult_21_n743), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n744), .ZN(p6_mult_21_n377) );
  XNOR2_X1 p6_mult_21_U561 ( .A(B0[2]), .B(reg1_reg[7]), .ZN(p6_mult_21_n744)
         );
  OAI22_X1 p6_mult_21_U490 ( .A1(p6_mult_21_n696), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n697), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n414) );
  XNOR2_X1 p6_mult_21_U493 ( .A(B0[8]), .B(reg1_reg[1]), .ZN(p6_mult_21_n697)
         );
  NOR2_X1 p6_mult_21_U582 ( .A1(p6_mult_21_n722), .A2(p6_mult_21_n757), .ZN(
        p6_mult_21_n365) );
  XNOR2_X1 p6_mult_21_U541 ( .A(B0[4]), .B(reg1_reg[5]), .ZN(p6_mult_21_n729)
         );
  OAI22_X1 p6_mult_21_U513 ( .A1(p6_mult_21_n711), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n712), .ZN(p6_mult_21_n402) );
  OAI22_X1 p6_mult_21_U488 ( .A1(p6_mult_21_n695), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n696), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n415) );
  XNOR2_X1 p6_mult_21_U491 ( .A(B0[7]), .B(reg1_reg[1]), .ZN(p6_mult_21_n696)
         );
  XNOR2_X1 p6_mult_21_U539 ( .A(B0[3]), .B(reg1_reg[5]), .ZN(p6_mult_21_n728)
         );
  XNOR2_X1 p6_mult_21_U559 ( .A(B0[1]), .B(reg1_reg[7]), .ZN(p6_mult_21_n743)
         );
  OAI22_X1 p6_mult_21_U511 ( .A1(p6_mult_21_n710), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n711), .ZN(p6_mult_21_n403) );
  NOR2_X1 p6_mult_21_U555 ( .A1(p6_mult_21_n722), .A2(p6_mult_21_n740), .ZN(
        p6_mult_21_n379) );
  OAI22_X1 p6_mult_21_U486 ( .A1(p6_mult_21_n694), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n695), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n416) );
  XNOR2_X1 p6_mult_21_U489 ( .A(B0[6]), .B(reg1_reg[1]), .ZN(p6_mult_21_n695)
         );
  XNOR2_X1 p6_mult_21_U537 ( .A(B0[2]), .B(reg1_reg[5]), .ZN(p6_mult_21_n727)
         );
  XNOR2_X1 p6_mult_21_U535 ( .A(B0[1]), .B(reg1_reg[5]), .ZN(p6_mult_21_n726)
         );
  XNOR2_X1 p6_mult_21_U533 ( .A(reg1_reg[5]), .B(B0[0]), .ZN(p6_mult_21_n724)
         );
  OAI21_X1 p6_mult_21_U659 ( .B1(p6_mult_21_n807), .B2(p6_mult_21_n725), .A(
        p6_mult_21_n808), .ZN(p6_mult_21_n321) );
  OAI22_X1 p6_mult_21_U484 ( .A1(p6_mult_21_n693), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n694), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n417) );
  XNOR2_X1 p6_mult_21_U487 ( .A(B0[5]), .B(reg1_reg[1]), .ZN(p6_mult_21_n694)
         );
  OAI22_X1 p6_mult_21_U509 ( .A1(p6_mult_21_n709), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n710), .ZN(p6_mult_21_n404) );
  OAI22_X1 p6_mult_21_U507 ( .A1(p6_mult_21_n708), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n709), .ZN(p6_mult_21_n405) );
  OAI22_X1 p6_mult_21_U482 ( .A1(p6_mult_21_n691), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n693), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n418) );
  XNOR2_X1 p6_mult_21_U485 ( .A(B0[4]), .B(reg1_reg[1]), .ZN(p6_mult_21_n693)
         );
  XNOR2_X1 p6_mult_21_U483 ( .A(B0[3]), .B(reg1_reg[1]), .ZN(p6_mult_21_n691)
         );
  NAND2_X1 p6_mult_21_U730 ( .A1(p6_mult_21_n842), .A2(p6_mult_21_n843), .ZN(
        p6_mult_21_n841) );
  NAND2_X1 p6_mult_21_U731 ( .A1(p6_mult_21_n837), .A2(p6_mult_21_n843), .ZN(
        p6_mult_21_n840) );
  OAI22_X1 p6_mult_21_U732 ( .A1(p6_mult_21_n844), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n689), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n843) );
  XNOR2_X1 p6_mult_21_U733 ( .A(B0[2]), .B(reg1_reg[1]), .ZN(p6_mult_21_n689)
         );
  NOR2_X1 p6_mult_21_U736 ( .A1(p6_mult_21_n704), .A2(B0[1]), .ZN(
        p6_mult_21_n842) );
  OAI22_X1 p6_mult_21_U496 ( .A1(p6_mult_21_n699), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n700), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n411) );
  XNOR2_X1 p6_mult_21_U497 ( .A(B0[10]), .B(reg1_reg[1]), .ZN(p6_mult_21_n699)
         );
  XNOR2_X1 p6_mult_21_U545 ( .A(B0[6]), .B(reg1_reg[5]), .ZN(p6_mult_21_n731)
         );
  OAI22_X1 p6_mult_21_U587 ( .A1(p6_mult_21_n761), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n762), .ZN(p6_mult_21_n362) );
  XNOR2_X1 p6_mult_21_U588 ( .A(B0[2]), .B(reg1_reg[9]), .ZN(p6_mult_21_n761)
         );
  XNOR2_X1 p6_mult_21_U547 ( .A(B0[7]), .B(reg1_reg[5]), .ZN(p6_mult_21_n732)
         );
  OAI22_X1 p6_mult_21_U566 ( .A1(p6_mult_21_n747), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n748), .ZN(p6_mult_21_n373) );
  XNOR2_X1 p6_mult_21_U567 ( .A(B0[5]), .B(reg1_reg[7]), .ZN(p6_mult_21_n747)
         );
  OAI22_X1 p6_mult_21_U523 ( .A1(p6_mult_21_n716), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n717), .ZN(p6_mult_21_n397) );
  OAI22_X1 p6_mult_21_U612 ( .A1(p6_mult_21_n777), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n778), .ZN(p6_mult_21_n349) );
  XNOR2_X1 p6_mult_21_U613 ( .A(B0[1]), .B(reg1_reg[11]), .ZN(p6_mult_21_n777)
         );
  OAI22_X1 p6_mult_21_U498 ( .A1(p6_mult_21_n700), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n701), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n410) );
  XNOR2_X1 p6_mult_21_U499 ( .A(B0[11]), .B(reg1_reg[1]), .ZN(p6_mult_21_n700)
         );
  NOR2_X1 p6_mult_21_U633 ( .A1(p6_mult_21_n722), .A2(p6_mult_21_n791), .ZN(
        p6_mult_21_n337) );
  OAI22_X1 p6_mult_21_U589 ( .A1(p6_mult_21_n762), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n763), .ZN(p6_mult_21_n361) );
  XNOR2_X1 p6_mult_21_U590 ( .A(B0[3]), .B(reg1_reg[9]), .ZN(p6_mult_21_n762)
         );
  OAI22_X1 p6_mult_21_U591 ( .A1(p6_mult_21_n763), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n764), .ZN(p6_mult_21_n360) );
  XNOR2_X1 p6_mult_21_U592 ( .A(B0[4]), .B(reg1_reg[9]), .ZN(p6_mult_21_n763)
         );
  XNOR2_X1 p6_mult_21_U549 ( .A(B0[8]), .B(reg1_reg[5]), .ZN(p6_mult_21_n733)
         );
  OAI22_X1 p6_mult_21_U614 ( .A1(p6_mult_21_n778), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n779), .ZN(p6_mult_21_n348) );
  XNOR2_X1 p6_mult_21_U615 ( .A(B0[2]), .B(reg1_reg[11]), .ZN(p6_mult_21_n778)
         );
  XNOR2_X1 p6_mult_21_U669 ( .A(p6_mult_21_n817), .B(p6_mult_21_n818), .ZN(
        p6_mult_21_n244) );
  OAI22_X1 p6_mult_21_U525 ( .A1(p6_mult_21_n717), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n718), .ZN(p6_mult_21_n396) );
  OAI22_X1 p6_mult_21_U568 ( .A1(p6_mult_21_n748), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n749), .ZN(p6_mult_21_n372) );
  XNOR2_X1 p6_mult_21_U569 ( .A(B0[6]), .B(reg1_reg[7]), .ZN(p6_mult_21_n748)
         );
  OAI22_X1 p6_mult_21_U500 ( .A1(p6_mult_21_n701), .A2(p6_mult_21_n690), .B1(
        p6_mult_21_n702), .B2(p6_mult_21_n692), .ZN(p6_mult_21_n409) );
  XNOR2_X1 p6_mult_21_U501 ( .A(B0[12]), .B(reg1_reg[1]), .ZN(p6_mult_21_n701)
         );
  OAI22_X1 p6_mult_21_U634 ( .A1(p6_mult_21_n792), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n794), .ZN(p6_mult_21_n336) );
  XNOR2_X1 p6_mult_21_U635 ( .A(reg1_reg[13]), .B(B0[0]), .ZN(p6_mult_21_n792)
         );
  OAI21_X1 p6_mult_21_U667 ( .B1(p6_mult_21_n815), .B2(p6_mult_21_n793), .A(
        p6_mult_21_n816), .ZN(p6_mult_21_n317) );
  OAI22_X1 p6_mult_21_U570 ( .A1(p6_mult_21_n749), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n750), .ZN(p6_mult_21_n371) );
  XNOR2_X1 p6_mult_21_U571 ( .A(B0[7]), .B(reg1_reg[7]), .ZN(p6_mult_21_n749)
         );
  OAI22_X1 p6_mult_21_U636 ( .A1(p6_mult_21_n794), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n795), .ZN(p6_mult_21_n335) );
  XNOR2_X1 p6_mult_21_U637 ( .A(B0[1]), .B(reg1_reg[13]), .ZN(p6_mult_21_n794)
         );
  XNOR2_X1 p6_mult_21_U673 ( .A(B0[9]), .B(reg1_reg[5]), .ZN(p6_mult_21_n734)
         );
  OAI22_X1 p6_mult_21_U674 ( .A1(p6_mult_21_n779), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n780), .ZN(p6_mult_21_n817) );
  XNOR2_X1 p6_mult_21_U676 ( .A(B0[3]), .B(reg1_reg[11]), .ZN(p6_mult_21_n779)
         );
  AOI21_X1 p6_mult_21_U503 ( .B1(p6_mult_21_n690), .B2(p6_mult_21_n692), .A(
        p6_mult_21_n702), .ZN(p6_mult_21_n703) );
  NAND2_X1 p6_mult_21_U734 ( .A1(reg1_reg[1]), .A2(p6_mult_21_n692), .ZN(
        p6_mult_21_n690) );
  OAI22_X1 p6_mult_21_U593 ( .A1(p6_mult_21_n764), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n765), .ZN(p6_mult_21_n359) );
  XNOR2_X1 p6_mult_21_U594 ( .A(B0[5]), .B(reg1_reg[9]), .ZN(p6_mult_21_n764)
         );
  OAI22_X1 p6_mult_21_U527 ( .A1(p6_mult_21_n718), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n719), .ZN(p6_mult_21_n395) );
  AOI21_X1 p6_mult_21_U530 ( .B1(p6_mult_21_n706), .B2(p6_mult_21_n707), .A(
        p6_mult_21_n721), .ZN(p6_mult_21_n720) );
  OAI22_X1 p6_mult_21_U640 ( .A1(p6_mult_21_n796), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n797), .ZN(p6_mult_21_n333) );
  OAI22_X1 p6_mult_21_U599 ( .A1(p6_mult_21_n767), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n768), .ZN(p6_mult_21_n356) );
  OAI22_X1 p6_mult_21_U642 ( .A1(p6_mult_21_n797), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n798), .ZN(p6_mult_21_n332) );
  XNOR2_X1 p6_mult_21_U643 ( .A(B0[4]), .B(reg1_reg[13]), .ZN(p6_mult_21_n797)
         );
  OAI22_X1 p6_mult_21_U595 ( .A1(p6_mult_21_n765), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n766), .ZN(p6_mult_21_n358) );
  XNOR2_X1 p6_mult_21_U596 ( .A(B0[6]), .B(reg1_reg[9]), .ZN(p6_mult_21_n765)
         );
  OAI22_X1 p6_mult_21_U572 ( .A1(p6_mult_21_n750), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n751), .ZN(p6_mult_21_n370) );
  XNOR2_X1 p6_mult_21_U573 ( .A(B0[8]), .B(reg1_reg[7]), .ZN(p6_mult_21_n750)
         );
  OAI22_X1 p6_mult_21_U638 ( .A1(p6_mult_21_n795), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n796), .ZN(p6_mult_21_n334) );
  XNOR2_X1 p6_mult_21_U641 ( .A(B0[3]), .B(reg1_reg[13]), .ZN(p6_mult_21_n796)
         );
  XNOR2_X1 p6_mult_21_U639 ( .A(B0[2]), .B(reg1_reg[13]), .ZN(p6_mult_21_n795)
         );
  OAI22_X1 p6_mult_21_U574 ( .A1(p6_mult_21_n751), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n752), .ZN(p6_mult_21_n369) );
  XNOR2_X1 p6_mult_21_U575 ( .A(B0[9]), .B(reg1_reg[7]), .ZN(p6_mult_21_n751)
         );
  OAI22_X1 p6_mult_21_U678 ( .A1(p6_mult_21_n719), .A2(p6_mult_21_n706), .B1(
        p6_mult_21_n707), .B2(p6_mult_21_n721), .ZN(p6_mult_21_n231) );
  XNOR2_X1 p6_mult_21_U725 ( .A(p6_mult_21_n820), .B(reg1_reg[2]), .ZN(
        p6_mult_21_n838) );
  OAI22_X1 p6_mult_21_U616 ( .A1(p6_mult_21_n780), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n781), .ZN(p6_mult_21_n346) );
  XNOR2_X1 p6_mult_21_U675 ( .A(B0[4]), .B(reg1_reg[11]), .ZN(p6_mult_21_n780)
         );
  XNOR2_X1 p6_mult_21_U672 ( .A(B0[10]), .B(reg1_reg[5]), .ZN(p6_mult_21_n735)
         );
  OAI22_X1 p6_mult_21_U597 ( .A1(p6_mult_21_n766), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n767), .ZN(p6_mult_21_n357) );
  XNOR2_X1 p6_mult_21_U600 ( .A(B0[8]), .B(reg1_reg[9]), .ZN(p6_mult_21_n767)
         );
  XNOR2_X1 p6_mult_21_U598 ( .A(B0[7]), .B(reg1_reg[9]), .ZN(p6_mult_21_n766)
         );
  XNOR2_X1 p6_mult_21_U552 ( .A(B0[11]), .B(reg1_reg[5]), .ZN(p6_mult_21_n736)
         );
  OAI22_X1 p6_mult_21_U617 ( .A1(p6_mult_21_n781), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n782), .ZN(p6_mult_21_n345) );
  XNOR2_X1 p6_mult_21_U618 ( .A(B0[5]), .B(reg1_reg[11]), .ZN(p6_mult_21_n781)
         );
  OAI22_X1 p6_mult_21_U619 ( .A1(p6_mult_21_n782), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n783), .ZN(p6_mult_21_n344) );
  XNOR2_X1 p6_mult_21_U620 ( .A(B0[6]), .B(reg1_reg[11]), .ZN(p6_mult_21_n782)
         );
  OAI22_X1 p6_mult_21_U576 ( .A1(p6_mult_21_n752), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n753), .ZN(p6_mult_21_n368) );
  XNOR2_X1 p6_mult_21_U577 ( .A(B0[10]), .B(reg1_reg[7]), .ZN(p6_mult_21_n752)
         );
  OAI22_X1 p6_mult_21_U578 ( .A1(p6_mult_21_n753), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n754), .ZN(p6_mult_21_n367) );
  XNOR2_X1 p6_mult_21_U579 ( .A(B0[11]), .B(reg1_reg[7]), .ZN(p6_mult_21_n753)
         );
  OAI22_X1 p6_mult_21_U621 ( .A1(p6_mult_21_n783), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n784), .ZN(p6_mult_21_n343) );
  XNOR2_X1 p6_mult_21_U622 ( .A(B0[7]), .B(reg1_reg[11]), .ZN(p6_mult_21_n783)
         );
  OAI22_X1 p6_mult_21_U601 ( .A1(p6_mult_21_n768), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n769), .ZN(p6_mult_21_n355) );
  XNOR2_X1 p6_mult_21_U602 ( .A(B0[9]), .B(reg1_reg[9]), .ZN(p6_mult_21_n768)
         );
  OAI22_X1 p6_mult_21_U603 ( .A1(p6_mult_21_n769), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n770), .ZN(p6_mult_21_n354) );
  XNOR2_X1 p6_mult_21_U604 ( .A(B0[10]), .B(reg1_reg[9]), .ZN(p6_mult_21_n769)
         );
  OAI22_X1 p6_mult_21_U644 ( .A1(p6_mult_21_n798), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n799), .ZN(p6_mult_21_n331) );
  XNOR2_X1 p6_mult_21_U645 ( .A(B0[5]), .B(reg1_reg[13]), .ZN(p6_mult_21_n798)
         );
  XNOR2_X1 p6_mult_21_U683 ( .A(B0[13]), .B(reg1_reg[5]), .ZN(p6_mult_21_n739)
         );
  XNOR2_X1 p6_mult_21_U684 ( .A(p6_mult_21_n807), .B(reg1_reg[4]), .ZN(
        p6_mult_21_n819) );
  XNOR2_X1 p6_mult_21_U685 ( .A(B0[12]), .B(reg1_reg[5]), .ZN(p6_mult_21_n737)
         );
  OAI22_X1 p6_mult_21_U623 ( .A1(p6_mult_21_n784), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n785), .ZN(p6_mult_21_n342) );
  XNOR2_X1 p6_mult_21_U624 ( .A(B0[8]), .B(reg1_reg[11]), .ZN(p6_mult_21_n784)
         );
  OAI22_X1 p6_mult_21_U646 ( .A1(p6_mult_21_n799), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n800), .ZN(p6_mult_21_n330) );
  XNOR2_X1 p6_mult_21_U647 ( .A(B0[6]), .B(reg1_reg[13]), .ZN(p6_mult_21_n799)
         );
  OAI22_X1 p6_mult_21_U605 ( .A1(p6_mult_21_n770), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n771), .ZN(p6_mult_21_n353) );
  XNOR2_X1 p6_mult_21_U606 ( .A(B0[11]), .B(reg1_reg[9]), .ZN(p6_mult_21_n770)
         );
  OAI22_X1 p6_mult_21_U625 ( .A1(p6_mult_21_n785), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n786), .ZN(p6_mult_21_n341) );
  XNOR2_X1 p6_mult_21_U626 ( .A(B0[9]), .B(reg1_reg[11]), .ZN(p6_mult_21_n785)
         );
  AOI21_X1 p6_mult_21_U581 ( .B1(p6_mult_21_n742), .B2(p6_mult_21_n740), .A(
        p6_mult_21_n756), .ZN(p6_mult_21_n755) );
  OAI22_X1 p6_mult_21_U648 ( .A1(p6_mult_21_n800), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n801), .ZN(p6_mult_21_n329) );
  XNOR2_X1 p6_mult_21_U649 ( .A(B0[7]), .B(reg1_reg[13]), .ZN(p6_mult_21_n800)
         );
  OAI22_X1 p6_mult_21_U687 ( .A1(p6_mult_21_n754), .A2(p6_mult_21_n742), .B1(
        p6_mult_21_n740), .B2(p6_mult_21_n756), .ZN(p6_mult_21_n191) );
  XNOR2_X1 p6_mult_21_U688 ( .A(B0[13]), .B(reg1_reg[7]), .ZN(p6_mult_21_n756)
         );
  XNOR2_X1 p6_mult_21_U690 ( .A(p6_mult_21_n809), .B(reg1_reg[6]), .ZN(
        p6_mult_21_n821) );
  XNOR2_X1 p6_mult_21_U692 ( .A(B0[12]), .B(reg1_reg[7]), .ZN(p6_mult_21_n754)
         );
  OAI22_X1 p6_mult_21_U629 ( .A1(p6_mult_21_n787), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n788), .ZN(p6_mult_21_n339) );
  OAI22_X1 p6_mult_21_U627 ( .A1(p6_mult_21_n786), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n787), .ZN(p6_mult_21_n340) );
  XNOR2_X1 p6_mult_21_U630 ( .A(B0[11]), .B(reg1_reg[11]), .ZN(p6_mult_21_n787) );
  XNOR2_X1 p6_mult_21_U628 ( .A(B0[10]), .B(reg1_reg[11]), .ZN(p6_mult_21_n786) );
  OAI22_X1 p6_mult_21_U650 ( .A1(p6_mult_21_n801), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n802), .ZN(p6_mult_21_n328) );
  XNOR2_X1 p6_mult_21_U651 ( .A(B0[8]), .B(reg1_reg[13]), .ZN(p6_mult_21_n801)
         );
  AOI21_X1 p6_mult_21_U608 ( .B1(p6_mult_21_n759), .B2(p6_mult_21_n757), .A(
        p6_mult_21_n773), .ZN(p6_mult_21_n772) );
  OAI22_X1 p6_mult_21_U694 ( .A1(p6_mult_21_n771), .A2(p6_mult_21_n759), .B1(
        p6_mult_21_n757), .B2(p6_mult_21_n773), .ZN(p6_mult_21_n177) );
  XNOR2_X1 p6_mult_21_U695 ( .A(B0[13]), .B(reg1_reg[9]), .ZN(p6_mult_21_n773)
         );
  XNOR2_X1 p6_mult_21_U697 ( .A(p6_mult_21_n811), .B(reg1_reg[8]), .ZN(
        p6_mult_21_n822) );
  XNOR2_X1 p6_mult_21_U699 ( .A(B0[12]), .B(reg1_reg[9]), .ZN(p6_mult_21_n771)
         );
  OAI22_X1 p6_mult_21_U652 ( .A1(p6_mult_21_n802), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n803), .ZN(p6_mult_21_n327) );
  XNOR2_X1 p6_mult_21_U653 ( .A(B0[9]), .B(reg1_reg[13]), .ZN(p6_mult_21_n802)
         );
  OAI22_X1 p6_mult_21_U654 ( .A1(p6_mult_21_n803), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n804), .ZN(p6_mult_21_n326) );
  XNOR2_X1 p6_mult_21_U655 ( .A(B0[10]), .B(reg1_reg[13]), .ZN(p6_mult_21_n803) );
  AOI22_X1 p6_mult_21_U707 ( .A1(p6_mult_21_n806), .A2(p6_mult_21_n686), .B1(
        p6_mult_21_n687), .B2(p6_mult_21_n688), .ZN(p6_mult_21_n162) );
  XNOR2_X1 p6_mult_21_U708 ( .A(B0[13]), .B(p6_mult_21_n815), .ZN(
        p6_mult_21_n688) );
  AOI21_X1 p6_mult_21_U632 ( .B1(p6_mult_21_n776), .B2(p6_mult_21_n774), .A(
        p6_mult_21_n790), .ZN(p6_mult_21_n789) );
  OAI22_X1 p6_mult_21_U701 ( .A1(p6_mult_21_n788), .A2(p6_mult_21_n776), .B1(
        p6_mult_21_n774), .B2(p6_mult_21_n790), .ZN(p6_mult_21_n167) );
  XNOR2_X1 p6_mult_21_U702 ( .A(B0[13]), .B(reg1_reg[11]), .ZN(p6_mult_21_n790) );
  XNOR2_X1 p6_mult_21_U704 ( .A(p6_mult_21_n813), .B(reg1_reg[10]), .ZN(
        p6_mult_21_n823) );
  XNOR2_X1 p6_mult_21_U706 ( .A(B0[12]), .B(reg1_reg[11]), .ZN(p6_mult_21_n788) );
  OAI22_X1 p6_mult_21_U656 ( .A1(p6_mult_21_n804), .A2(p6_mult_21_n793), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n805), .ZN(p6_mult_21_n325) );
  XNOR2_X1 p6_mult_21_U712 ( .A(p6_mult_21_n815), .B(reg1_reg[12]), .ZN(
        p6_mult_21_n824) );
  XNOR2_X1 p6_mult_21_U658 ( .A(B0[11]), .B(reg1_reg[13]), .ZN(p6_mult_21_n804) );
  XOR2_X1 p6_mult_21_U738 ( .A(reg1_reg[2]), .B(reg1_reg[1]), .Z(
        p6_mult_21_n837) );
  MUX2_X1 p6_mult_21_U728 ( .A(p6_mult_21_n840), .B(p6_mult_21_n841), .S(
        p6_mult_21_n722), .Z(p6_mult_21_n839) );
  XOR2_X1 p6_mult_21_U715 ( .A(B0[12]), .B(reg1_reg[13]), .Z(p6_mult_21_n806)
         );
  NAND3_X1 p6_mult_21_U668 ( .A1(p6_mult_21_n687), .A2(p6_mult_21_n722), .A3(
        reg1_reg[13]), .ZN(p6_mult_21_n816) );
  XOR2_X1 p6_mult_21_U504 ( .A(B0[13]), .B(p6_mult_21_n704), .Z(
        p6_mult_21_n702) );
  NAND3_X1 p6_mult_21_U465 ( .A1(p6_mult_21_n672), .A2(p6_mult_21_n673), .A3(
        p6_mult_21_n674), .ZN(p6_mult_21_n148) );
  XOR2_X1 p6_mult_21_U461 ( .A(p6_mult_21_n640), .B(p6_mult_21_n671), .Z(
        temp1[0]) );
  XOR2_X1 p6_mult_21_U460 ( .A(p6_mult_21_n246), .B(p6_mult_21_n257), .Z(
        p6_mult_21_n671) );
  XOR2_X1 p6_mult_21_U455 ( .A(p6_mult_21_n148), .B(p6_mult_21_n667), .Z(
        temp1[1]) );
  XOR2_X1 p6_mult_21_U454 ( .A(p6_mult_21_n234), .B(p6_mult_21_n245), .Z(
        p6_mult_21_n667) );
  XOR2_X1 p6_mult_21_U435 ( .A(p6_mult_21_n141), .B(p6_mult_21_n651), .Z(
        temp1[8]) );
  XOR2_X1 p6_mult_21_U434 ( .A(p6_mult_21_n179), .B(p6_mult_21_n174), .Z(
        p6_mult_21_n651) );
  XOR2_X1 p6_mult_21_U429 ( .A(p6_mult_21_n142), .B(p6_mult_21_n647), .Z(
        temp1[7]) );
  XOR2_X1 p6_mult_21_U428 ( .A(p6_mult_21_n180), .B(p6_mult_21_n185), .Z(
        p6_mult_21_n647) );
  NAND3_X1 p6_mult_21_U409 ( .A1(p6_mult_21_n641), .A2(p6_mult_21_n642), .A3(
        p6_mult_21_n643), .ZN(p6_mult_21_n635) );
  FA_X1 p6_mult_21_U144 ( .A(p6_mult_21_n418), .B(p6_mult_21_n393), .CI(
        p6_mult_21_n405), .CO(p6_mult_21_n313), .S(p6_mult_21_n314) );
  HA_X1 p6_mult_21_U143 ( .A(p6_mult_21_n321), .B(p6_mult_21_n392), .CO(
        p6_mult_21_n311), .S(p6_mult_21_n312) );
  FA_X1 p6_mult_21_U141 ( .A(p6_mult_21_n416), .B(p6_mult_21_n379), .CI(
        p6_mult_21_n403), .CO(p6_mult_21_n307), .S(p6_mult_21_n308) );
  FA_X1 p6_mult_21_U138 ( .A(p6_mult_21_n390), .B(p6_mult_21_n415), .CI(
        p6_mult_21_n402), .CO(p6_mult_21_n301), .S(p6_mult_21_n302) );
  FA_X1 p6_mult_21_U137 ( .A(p6_mult_21_n307), .B(p6_mult_21_n304), .CI(
        p6_mult_21_n302), .CO(p6_mult_21_n299), .S(p6_mult_21_n300) );
  FA_X1 p6_mult_21_U136 ( .A(p6_mult_21_n389), .B(p6_mult_21_n365), .CI(
        p6_mult_21_n414), .CO(p6_mult_21_n297), .S(p6_mult_21_n298) );
  FA_X1 p6_mult_21_U135 ( .A(p6_mult_21_n377), .B(p6_mult_21_n401), .CI(
        p6_mult_21_n303), .CO(p6_mult_21_n295), .S(p6_mult_21_n296) );
  FA_X1 p6_mult_21_U134 ( .A(p6_mult_21_n298), .B(p6_mult_21_n301), .CI(
        p6_mult_21_n296), .CO(p6_mult_21_n293), .S(p6_mult_21_n294) );
  FA_X1 p6_mult_21_U132 ( .A(p6_mult_21_n376), .B(p6_mult_21_n388), .CI(
        p6_mult_21_n400), .CO(p6_mult_21_n289), .S(p6_mult_21_n290) );
  FA_X1 p6_mult_21_U131 ( .A(p6_mult_21_n292), .B(p6_mult_21_n413), .CI(
        p6_mult_21_n297), .CO(p6_mult_21_n287), .S(p6_mult_21_n288) );
  FA_X1 p6_mult_21_U130 ( .A(p6_mult_21_n290), .B(p6_mult_21_n295), .CI(
        p6_mult_21_n288), .CO(p6_mult_21_n285), .S(p6_mult_21_n286) );
  FA_X1 p6_mult_21_U129 ( .A(p6_mult_21_n375), .B(p6_mult_21_n351), .CI(
        p6_mult_21_n412), .CO(p6_mult_21_n283), .S(p6_mult_21_n284) );
  FA_X1 p6_mult_21_U128 ( .A(p6_mult_21_n363), .B(p6_mult_21_n399), .CI(
        p6_mult_21_n387), .CO(p6_mult_21_n281), .S(p6_mult_21_n282) );
  FA_X1 p6_mult_21_U127 ( .A(p6_mult_21_n289), .B(p6_mult_21_n291), .CI(
        p6_mult_21_n284), .CO(p6_mult_21_n279), .S(p6_mult_21_n280) );
  FA_X1 p6_mult_21_U126 ( .A(p6_mult_21_n287), .B(p6_mult_21_n282), .CI(
        p6_mult_21_n280), .CO(p6_mult_21_n277), .S(p6_mult_21_n278) );
  FA_X1 p6_mult_21_U124 ( .A(p6_mult_21_n362), .B(p6_mult_21_n386), .CI(
        p6_mult_21_n411), .CO(p6_mult_21_n273), .S(p6_mult_21_n274) );
  FA_X1 p6_mult_21_U123 ( .A(p6_mult_21_n374), .B(p6_mult_21_n398), .CI(
        p6_mult_21_n276), .CO(p6_mult_21_n271), .S(p6_mult_21_n272) );
  FA_X1 p6_mult_21_U122 ( .A(p6_mult_21_n281), .B(p6_mult_21_n283), .CI(
        p6_mult_21_n274), .CO(p6_mult_21_n269), .S(p6_mult_21_n270) );
  FA_X1 p6_mult_21_U121 ( .A(p6_mult_21_n279), .B(p6_mult_21_n272), .CI(
        p6_mult_21_n270), .CO(p6_mult_21_n267), .S(p6_mult_21_n268) );
  FA_X1 p6_mult_21_U120 ( .A(p6_mult_21_n361), .B(p6_mult_21_n337), .CI(
        p6_mult_21_n410), .CO(p6_mult_21_n265), .S(p6_mult_21_n266) );
  FA_X1 p6_mult_21_U109 ( .A(p6_mult_21_n349), .B(p6_mult_21_n397), .CI(
        p6_mult_21_n373), .CO(p6_mult_21_n263), .S(p6_mult_21_n264) );
  FA_X1 p6_mult_21_U108 ( .A(p6_mult_21_n275), .B(p6_mult_21_n385), .CI(
        p6_mult_21_n273), .CO(p6_mult_21_n261), .S(p6_mult_21_n262) );
  FA_X1 p6_mult_21_U107 ( .A(p6_mult_21_n264), .B(p6_mult_21_n266), .CI(
        p6_mult_21_n271), .CO(p6_mult_21_n259), .S(p6_mult_21_n260) );
  FA_X1 p6_mult_21_U106 ( .A(p6_mult_21_n262), .B(p6_mult_21_n269), .CI(
        p6_mult_21_n260), .CO(p6_mult_21_n257), .S(p6_mult_21_n258) );
  HA_X1 p6_mult_21_U105 ( .A(p6_mult_21_n317), .B(p6_mult_21_n336), .CO(
        p6_mult_21_n255), .S(p6_mult_21_n256) );
  FA_X1 p6_mult_21_U104 ( .A(p6_mult_21_n409), .B(p6_mult_21_n372), .CI(
        p6_mult_21_n396), .CO(p6_mult_21_n253), .S(p6_mult_21_n254) );
  FA_X1 p6_mult_21_U103 ( .A(p6_mult_21_n348), .B(p6_mult_21_n384), .CI(
        p6_mult_21_n360), .CO(p6_mult_21_n251), .S(p6_mult_21_n252) );
  FA_X1 p6_mult_21_U102 ( .A(p6_mult_21_n265), .B(p6_mult_21_n256), .CI(
        p6_mult_21_n263), .CO(p6_mult_21_n249), .S(p6_mult_21_n250) );
  FA_X1 p6_mult_21_U101 ( .A(p6_mult_21_n254), .B(p6_mult_21_n252), .CI(
        p6_mult_21_n261), .CO(p6_mult_21_n247), .S(p6_mult_21_n248) );
  FA_X1 p6_mult_21_U100 ( .A(p6_mult_21_n259), .B(p6_mult_21_n250), .CI(
        p6_mult_21_n248), .CO(p6_mult_21_n245), .S(p6_mult_21_n246) );
  FA_X1 p6_mult_21_U97 ( .A(p6_mult_21_n395), .B(p6_mult_21_n359), .CI(
        p6_mult_21_n408), .CO(p6_mult_21_n241), .S(p6_mult_21_n242) );
  FA_X1 p6_mult_21_U96 ( .A(p6_mult_21_n335), .B(p6_mult_21_n371), .CI(
        p6_mult_21_n255), .CO(p6_mult_21_n239), .S(p6_mult_21_n240) );
  FA_X1 p6_mult_21_U95 ( .A(p6_mult_21_n253), .B(p6_mult_21_n244), .CI(
        p6_mult_21_n251), .CO(p6_mult_21_n237), .S(p6_mult_21_n238) );
  FA_X1 p6_mult_21_U94 ( .A(p6_mult_21_n240), .B(p6_mult_21_n242), .CI(
        p6_mult_21_n249), .CO(p6_mult_21_n235), .S(p6_mult_21_n236) );
  FA_X1 p6_mult_21_U93 ( .A(p6_mult_21_n247), .B(p6_mult_21_n238), .CI(
        p6_mult_21_n236), .CO(p6_mult_21_n233), .S(p6_mult_21_n234) );
  FA_X1 p6_mult_21_U91 ( .A(p6_mult_21_n382), .B(p6_mult_21_n346), .CI(
        p6_mult_21_n232), .CO(p6_mult_21_n229), .S(p6_mult_21_n230) );
  FA_X1 p6_mult_21_U90 ( .A(p6_mult_21_n334), .B(p6_mult_21_n370), .CI(
        p6_mult_21_n358), .CO(p6_mult_21_n227), .S(p6_mult_21_n228) );
  FA_X1 p6_mult_21_U89 ( .A(p6_mult_21_n241), .B(p6_mult_21_n243), .CI(
        p6_mult_21_n239), .CO(p6_mult_21_n225), .S(p6_mult_21_n226) );
  FA_X1 p6_mult_21_U88 ( .A(p6_mult_21_n230), .B(p6_mult_21_n228), .CI(
        p6_mult_21_n237), .CO(p6_mult_21_n223), .S(p6_mult_21_n224) );
  FA_X1 p6_mult_21_U87 ( .A(p6_mult_21_n235), .B(p6_mult_21_n226), .CI(
        p6_mult_21_n224), .CO(p6_mult_21_n221), .S(p6_mult_21_n222) );
  FA_X1 p6_mult_21_U86 ( .A(p6_mult_21_n231), .B(p6_mult_21_n333), .CI(
        p6_mult_21_n394), .CO(p6_mult_21_n219), .S(p6_mult_21_n220) );
  FA_X1 p6_mult_21_U85 ( .A(p6_mult_21_n345), .B(p6_mult_21_n381), .CI(
        p6_mult_21_n357), .CO(p6_mult_21_n217), .S(p6_mult_21_n218) );
  FA_X1 p6_mult_21_U84 ( .A(p6_mult_21_n229), .B(p6_mult_21_n369), .CI(
        p6_mult_21_n227), .CO(p6_mult_21_n215), .S(p6_mult_21_n216) );
  FA_X1 p6_mult_21_U83 ( .A(p6_mult_21_n220), .B(p6_mult_21_n218), .CI(
        p6_mult_21_n225), .CO(p6_mult_21_n213), .S(p6_mult_21_n214) );
  FA_X1 p6_mult_21_U82 ( .A(p6_mult_21_n223), .B(p6_mult_21_n216), .CI(
        p6_mult_21_n214), .CO(p6_mult_21_n211), .S(p6_mult_21_n212) );
  FA_X1 p6_mult_21_U80 ( .A(p6_mult_21_n368), .B(p6_mult_21_n344), .CI(
        p6_mult_21_n210), .CO(p6_mult_21_n207), .S(p6_mult_21_n208) );
  FA_X1 p6_mult_21_U79 ( .A(p6_mult_21_n332), .B(p6_mult_21_n356), .CI(
        p6_mult_21_n219), .CO(p6_mult_21_n205), .S(p6_mult_21_n206) );
  FA_X1 p6_mult_21_U78 ( .A(p6_mult_21_n208), .B(p6_mult_21_n217), .CI(
        p6_mult_21_n215), .CO(p6_mult_21_n203), .S(p6_mult_21_n204) );
  FA_X1 p6_mult_21_U77 ( .A(p6_mult_21_n213), .B(p6_mult_21_n206), .CI(
        p6_mult_21_n204), .CO(p6_mult_21_n201), .S(p6_mult_21_n202) );
  FA_X1 p6_mult_21_U76 ( .A(p6_mult_21_n209), .B(p6_mult_21_n331), .CI(
        p6_mult_21_n380), .CO(p6_mult_21_n199), .S(p6_mult_21_n200) );
  FA_X1 p6_mult_21_U75 ( .A(p6_mult_21_n355), .B(p6_mult_21_n343), .CI(
        p6_mult_21_n367), .CO(p6_mult_21_n197), .S(p6_mult_21_n198) );
  FA_X1 p6_mult_21_U74 ( .A(p6_mult_21_n198), .B(p6_mult_21_n207), .CI(
        p6_mult_21_n200), .CO(p6_mult_21_n195), .S(p6_mult_21_n196) );
  FA_X1 p6_mult_21_U73 ( .A(p6_mult_21_n203), .B(p6_mult_21_n205), .CI(
        p6_mult_21_n196), .CO(p6_mult_21_n193), .S(p6_mult_21_n194) );
  FA_X1 p6_mult_21_U71 ( .A(p6_mult_21_n330), .B(p6_mult_21_n342), .CI(
        p6_mult_21_n192), .CO(p6_mult_21_n189), .S(p6_mult_21_n190) );
  FA_X1 p6_mult_21_U70 ( .A(p6_mult_21_n199), .B(p6_mult_21_n354), .CI(
        p6_mult_21_n197), .CO(p6_mult_21_n187), .S(p6_mult_21_n188) );
  FA_X1 p6_mult_21_U69 ( .A(p6_mult_21_n188), .B(p6_mult_21_n190), .CI(
        p6_mult_21_n195), .CO(p6_mult_21_n185), .S(p6_mult_21_n186) );
  FA_X1 p6_mult_21_U68 ( .A(p6_mult_21_n191), .B(p6_mult_21_n329), .CI(
        p6_mult_21_n366), .CO(p6_mult_21_n183), .S(p6_mult_21_n184) );
  FA_X1 p6_mult_21_U67 ( .A(p6_mult_21_n341), .B(p6_mult_21_n353), .CI(
        p6_mult_21_n189), .CO(p6_mult_21_n181), .S(p6_mult_21_n182) );
  FA_X1 p6_mult_21_U66 ( .A(p6_mult_21_n187), .B(p6_mult_21_n184), .CI(
        p6_mult_21_n182), .CO(p6_mult_21_n179), .S(p6_mult_21_n180) );
  FA_X1 p6_mult_21_U64 ( .A(p6_mult_21_n328), .B(p6_mult_21_n340), .CI(
        p6_mult_21_n178), .CO(p6_mult_21_n175), .S(p6_mult_21_n176) );
  FA_X1 p6_mult_21_U63 ( .A(p6_mult_21_n176), .B(p6_mult_21_n183), .CI(
        p6_mult_21_n181), .CO(p6_mult_21_n173), .S(p6_mult_21_n174) );
  FA_X1 p6_mult_21_U62 ( .A(p6_mult_21_n327), .B(p6_mult_21_n177), .CI(
        p6_mult_21_n352), .CO(p6_mult_21_n171), .S(p6_mult_21_n172) );
  FA_X1 p6_mult_21_U61 ( .A(p6_mult_21_n175), .B(p6_mult_21_n339), .CI(
        p6_mult_21_n172), .CO(p6_mult_21_n169), .S(p6_mult_21_n170) );
  FA_X1 p6_mult_21_U59 ( .A(p6_mult_21_n168), .B(p6_mult_21_n326), .CI(
        p6_mult_21_n171), .CO(p6_mult_21_n165), .S(p6_mult_21_n166) );
  FA_X1 p6_mult_21_U58 ( .A(p6_mult_21_n325), .B(p6_mult_21_n167), .CI(
        p6_mult_21_n338), .CO(p6_mult_21_n163), .S(p6_mult_21_n164) );
  FA_X1 p6_mult_21_U42 ( .A(p6_mult_21_n222), .B(p6_mult_21_n233), .CI(
        p6_mult_21_n147), .CO(p6_mult_21_n146), .S(temp1[2]) );
  FA_X1 p6_mult_21_U41 ( .A(p6_mult_21_n212), .B(p6_mult_21_n221), .CI(
        p6_mult_21_n146), .CO(p6_mult_21_n145), .S(temp1[3]) );
  FA_X1 p6_mult_21_U40 ( .A(p6_mult_21_n202), .B(p6_mult_21_n211), .CI(
        p6_mult_21_n145), .CO(p6_mult_21_n144), .S(temp1[4]) );
  FA_X1 p6_mult_21_U39 ( .A(p6_mult_21_n194), .B(p6_mult_21_n201), .CI(
        p6_mult_21_n144), .CO(p6_mult_21_n143), .S(temp1[5]) );
  FA_X1 p6_mult_21_U38 ( .A(p6_mult_21_n186), .B(p6_mult_21_n193), .CI(
        p6_mult_21_n143), .CO(p6_mult_21_n142), .S(temp1[6]) );
  FA_X1 p6_mult_21_U20 ( .A(p6_mult_21_n170), .B(p6_mult_21_n173), .CI(
        p6_mult_21_n140), .CO(p6_mult_21_n139), .S(temp1[9]) );
  FA_X1 p6_mult_21_U10 ( .A(p6_mult_21_n166), .B(p6_mult_21_n169), .CI(
        p6_mult_21_n139), .CO(p6_mult_21_n138), .S(temp1[10]) );
  FA_X1 p6_mult_21_U9 ( .A(p6_mult_21_n165), .B(p6_mult_21_n164), .CI(
        p6_mult_21_n138), .CO(p6_mult_21_n137), .S(temp1[11]) );
  FA_X1 p6_mult_21_U8 ( .A(p6_mult_21_n163), .B(p6_mult_21_n162), .CI(
        p6_mult_21_n137), .CO(p6_mult_21_n136), .S(temp1[12]) );
  INV_X1 p7_mult_21_U446 ( .A(p7_mult_21_n884), .ZN(p7_mult_21_n902) );
  INV_X1 p7_mult_21_U457 ( .A(p7_mult_21_n922), .ZN(p7_mult_21_n906) );
  INV_X1 p7_mult_21_U514 ( .A(p7_mult_21_n1008), .ZN(p7_mult_21_n1005) );
  INV_X1 p7_mult_21_U540 ( .A(p7_mult_21_n1000), .ZN(p7_mult_21_n1026) );
  INV_X1 p7_mult_21_U549 ( .A(p7_mult_21_n1061), .ZN(p7_mult_21_n1059) );
  INV_X1 p7_mult_21_U779 ( .A(p7_mult_21_n1361), .ZN(p7_mult_21_n1367) );
  INV_X1 p7_mult_21_U790 ( .A(p7_mult_21_n1372), .ZN(p7_mult_21_n1371) );
  INV_X1 p7_mult_21_U765 ( .A(p7_mult_21_n1352), .ZN(p7_mult_21_n1202) );
  INV_X1 p7_mult_21_U838 ( .A(p7_mult_21_n1396), .ZN(p7_mult_21_n1395) );
  INV_X1 p7_mult_21_U832 ( .A(p7_mult_21_n1393), .ZN(p7_mult_21_n1206) );
  INV_X1 p7_mult_21_U649 ( .A(p7_mult_21_n1211), .ZN(p7_mult_21_n1210) );
  INV_X1 p7_mult_21_U653 ( .A(p7_mult_21_n1221), .ZN(p7_mult_21_n1220) );
  AND2_X1 p7_mult_21_U683 ( .A1(p7_mult_21_n1277), .A2(p7_mult_21_n1278), .ZN(
        p7_mult_21_n1232) );
  INV_X1 p7_mult_21_U691 ( .A(p7_mult_21_n1286), .ZN(p7_mult_21_n1250) );
  INV_X1 p7_mult_21_U770 ( .A(p7_mult_21_n1344), .ZN(p7_mult_21_n1355) );
  INV_X1 p7_mult_21_U723 ( .A(p7_mult_21_n1328), .ZN(p7_mult_21_n1326) );
  AND2_X1 p7_mult_21_U740 ( .A1(p7_mult_21_n1302), .A2(p7_mult_21_n1303), .ZN(
        p7_mult_21_n1298) );
  INV_X1 p7_mult_21_U748 ( .A(p7_mult_21_n1342), .ZN(p7_mult_21_n1341) );
  INV_X1 p7_mult_21_U868 ( .A(p7_mult_21_n1402), .ZN(p7_mult_21_n1390) );
  INV_X1 p7_mult_21_U749 ( .A(p7_mult_21_n1028), .ZN(p7_mult_21_n1089) );
  INV_X1 p7_mult_21_U573 ( .A(p7_mult_21_n1066), .ZN(p7_mult_21_n1092) );
  INV_X1 p7_mult_21_U577 ( .A(p7_mult_21_n1067), .ZN(p7_mult_21_n1098) );
  AND2_X1 p7_mult_21_U605 ( .A1(p7_mult_21_n1135), .A2(p7_mult_21_n1136), .ZN(
        p7_mult_21_n1103) );
  INV_X1 p7_mult_21_U629 ( .A(p7_mult_21_n1172), .ZN(p7_mult_21_n1171) );
  AND2_X1 p7_mult_21_U632 ( .A1(p7_mult_21_n1177), .A2(p7_mult_21_n1178), .ZN(
        p7_mult_21_n1140) );
  INV_X1 p7_mult_21_U588 ( .A(p7_mult_21_n1090), .ZN(p7_mult_21_n1121) );
  INV_X1 p7_mult_21_U594 ( .A(p7_mult_21_n1091), .ZN(p7_mult_21_n1127) );
  INV_X1 p7_mult_21_U794 ( .A(p7_mult_21_n1376), .ZN(p7_mult_21_n1162) );
  INV_X1 p7_mult_21_U586 ( .A(p7_mult_21_n1119), .ZN(p7_mult_21_n1116) );
  INV_X1 p7_mult_21_U860 ( .A(p7_mult_21_n1096), .ZN(p7_mult_21_n1124) );
  INV_X1 p7_mult_21_U808 ( .A(p7_mult_21_n1289), .ZN(p7_mult_21_n1271) );
  INV_X1 p7_mult_21_U508 ( .A(p7_mult_21_n971), .ZN(p7_mult_21_n996) );
  INV_X1 p7_mult_21_U747 ( .A(p7_mult_21_n1029), .ZN(p7_mult_21_n1051) );
  INV_X1 p7_mult_21_U511 ( .A(p7_mult_21_n1001), .ZN(p7_mult_21_n999) );
  INV_X1 p7_mult_21_U847 ( .A(B1[5]), .ZN(p7_mult_21_n1068) );
  INV_X1 p7_mult_21_U852 ( .A(p7_mult_21_n957), .ZN(p7_mult_21_n1022) );
  INV_X1 p7_mult_21_U521 ( .A(p7_mult_21_n1020), .ZN(p7_mult_21_n1002) );
  INV_X1 p7_mult_21_U472 ( .A(p7_mult_21_n946), .ZN(p7_mult_21_n917) );
  INV_X1 p7_mult_21_U817 ( .A(B1[11]), .ZN(p7_mult_21_n904) );
  INV_X1 p7_mult_21_U880 ( .A(p7_mult_21_n920), .ZN(p7_mult_21_n943) );
  INV_X1 p7_mult_21_U885 ( .A(p7_mult_21_n919), .ZN(p7_mult_21_n970) );
  INV_X1 p7_mult_21_U864 ( .A(B1[10]), .ZN(p7_mult_21_n924) );
  INV_X1 p7_mult_21_U501 ( .A(p7_mult_21_n993), .ZN(p7_mult_21_n969) );
  INV_X1 p7_mult_21_U843 ( .A(p7_mult_21_n887), .ZN(p7_mult_21_n909) );
  AOI221_X1 p7_mult_21_U872 ( .B1(reg2_reg[10]), .B2(reg2_reg[11]), .C1(
        p7_mult_21_n1403), .C2(p7_mult_21_n911), .A(p7_mult_21_n886), .ZN(
        p7_mult_21_n887) );
  INV_X1 p7_mult_21_U859 ( .A(B1[9]), .ZN(p7_mult_21_n941) );
  INV_X1 p7_mult_21_U764 ( .A(p7_mult_21_n886), .ZN(p7_mult_21_n914) );
  INV_X1 p7_mult_21_U851 ( .A(B1[6]), .ZN(p7_mult_21_n1032) );
  INV_X1 p7_mult_21_U848 ( .A(p7_mult_21_n958), .ZN(p7_mult_21_n990) );
  INV_X1 p7_mult_21_U897 ( .A(B1[12]), .ZN(p7_mult_21_n885) );
  INV_X1 p7_mult_21_U480 ( .A(p7_mult_21_n960), .ZN(p7_mult_21_n952) );
  INV_X1 p7_mult_21_U814 ( .A(B1[7]), .ZN(p7_mult_21_n988) );
  INV_X1 p7_mult_21_U822 ( .A(p7_mult_21_n874), .ZN(p7_mult_21_n867) );
  INV_X1 p7_mult_21_U837 ( .A(B1[8]), .ZN(p7_mult_21_n962) );
  INV_X1 p7_mult_21_U557 ( .A(p7_mult_21_n883), .ZN(p7_mult_21_n866) );
  INV_X1 p7_mult_21_U811 ( .A(B1[13]), .ZN(p7_mult_21_n877) );
  AOI221_X1 p7_mult_21_U881 ( .B1(reg2_reg[8]), .B2(reg2_reg[9]), .C1(
        p7_mult_21_n1331), .C2(p7_mult_21_n945), .A(p7_mult_21_n919), .ZN(
        p7_mult_21_n920) );
  AOI22_X1 p7_mult_21_U886 ( .A1(reg2_reg[8]), .A2(reg2_reg[7]), .B1(
        p7_mult_21_n992), .B2(p7_mult_21_n1331), .ZN(p7_mult_21_n919) );
  AOI22_X1 p7_mult_21_U875 ( .A1(reg2_reg[9]), .A2(reg2_reg[10]), .B1(
        p7_mult_21_n1403), .B2(p7_mult_21_n945), .ZN(p7_mult_21_n886) );
  AOI22_X1 p7_mult_21_U891 ( .A1(reg2_reg[12]), .A2(p7_mult_21_n911), .B1(
        reg2_reg[11]), .B2(p7_mult_21_n1386), .ZN(p7_mult_21_n883) );
  XNOR2_X1 p7_mult_21_U612 ( .A(p7_mult_21_n1108), .B(p7_mult_21_n1110), .ZN(
        p7_mult_21_n1146) );
  XNOR2_X1 p7_mult_21_U637 ( .A(p7_mult_21_n1149), .B(p7_mult_21_n1182), .ZN(
        temp2[0]) );
  XNOR2_X1 p7_mult_21_U581 ( .A(p7_mult_21_n1075), .B(p7_mult_21_n1107), .ZN(
        temp2[2]) );
  XNOR2_X1 p7_mult_21_U561 ( .A(p7_mult_21_n1040), .B(p7_mult_21_n1041), .ZN(
        p7_mult_21_n1072) );
  XNOR2_X1 p7_mult_21_U533 ( .A(p7_mult_21_n1035), .B(p7_mult_21_n1039), .ZN(
        temp2[4]) );
  XNOR2_X1 p7_mult_21_U515 ( .A(p7_mult_21_n1009), .B(p7_mult_21_n981), .ZN(
        temp2[5]) );
  XNOR2_X1 p7_mult_21_U492 ( .A(p7_mult_21_n974), .B(p7_mult_21_n978), .ZN(
        temp2[6]) );
  XNOR2_X1 p7_mult_21_U478 ( .A(p7_mult_21_n954), .B(p7_mult_21_n934), .ZN(
        temp2[7]) );
  XNOR2_X1 p7_mult_21_U463 ( .A(p7_mult_21_n927), .B(p7_mult_21_n931), .ZN(
        temp2[8]) );
  XNOR2_X1 p7_mult_21_U452 ( .A(p7_mult_21_n912), .B(p7_mult_21_n897), .ZN(
        temp2[9]) );
  XNOR2_X1 p7_mult_21_U442 ( .A(p7_mult_21_n891), .B(p7_mult_21_n894), .ZN(
        temp2[10]) );
  OAI21_X1 p7_mult_21_U431 ( .B1(p7_mult_21_n873), .B2(p7_mult_21_n874), .A(
        p7_mult_21_n875), .ZN(p7_mult_21_n860) );
  NAND2_X1 p7_mult_21_U432 ( .A1(p7_mult_21_n868), .A2(p7_mult_21_n866), .ZN(
        p7_mult_21_n875) );
  AOI22_X1 p7_mult_21_U433 ( .A1(B1[13]), .A2(reg2_reg[13]), .B1(
        p7_mult_21_n876), .B2(p7_mult_21_n877), .ZN(p7_mult_21_n868) );
  AOI222_X1 p7_mult_21_U430 ( .A1(p7_mult_21_n870), .A2(p7_mult_21_n871), .B1(
        p7_mult_21_n870), .B2(p7_mult_21_n872), .C1(p7_mult_21_n871), .C2(
        p7_mult_21_n872), .ZN(p7_mult_21_n864) );
  AOI222_X1 p7_mult_21_U441 ( .A1(p7_mult_21_n892), .A2(p7_mult_21_n893), .B1(
        p7_mult_21_n892), .B2(p7_mult_21_n872), .C1(p7_mult_21_n893), .C2(
        p7_mult_21_n872), .ZN(p7_mult_21_n878) );
  OAI22_X1 p7_mult_21_U436 ( .A1(p7_mult_21_n883), .A2(p7_mult_21_n873), .B1(
        p7_mult_21_n874), .B2(p7_mult_21_n884), .ZN(p7_mult_21_n871) );
  AOI22_X1 p7_mult_21_U437 ( .A1(reg2_reg[13]), .A2(p7_mult_21_n885), .B1(
        B1[12]), .B2(p7_mult_21_n876), .ZN(p7_mult_21_n873) );
  OAI21_X1 p7_mult_21_U438 ( .B1(p7_mult_21_n886), .B2(n673), .A(
        p7_mult_21_n888), .ZN(p7_mult_21_n870) );
  AOI22_X1 p7_mult_21_U445 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n902), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n903), .ZN(p7_mult_21_n893) );
  AOI22_X1 p7_mult_21_U447 ( .A1(reg2_reg[13]), .A2(p7_mult_21_n904), .B1(
        B1[11]), .B2(p7_mult_21_n876), .ZN(p7_mult_21_n884) );
  AOI222_X1 p7_mult_21_U448 ( .A1(p7_mult_21_n905), .A2(p7_mult_21_n906), .B1(
        p7_mult_21_n905), .B2(p7_mult_21_n907), .C1(p7_mult_21_n906), .C2(
        p7_mult_21_n907), .ZN(p7_mult_21_n892) );
  OAI21_X1 p7_mult_21_U449 ( .B1(p7_mult_21_n908), .B2(p7_mult_21_n909), .A(
        p7_mult_21_n910), .ZN(p7_mult_21_n872) );
  NAND2_X1 p7_mult_21_U450 ( .A1(p7_mult_21_n886), .A2(p7_mult_21_n888), .ZN(
        p7_mult_21_n910) );
  AOI22_X1 p7_mult_21_U451 ( .A1(B1[13]), .A2(reg2_reg[11]), .B1(
        p7_mult_21_n911), .B2(p7_mult_21_n877), .ZN(p7_mult_21_n888) );
  OAI22_X1 p7_mult_21_U453 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n908), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n915), .ZN(p7_mult_21_n899) );
  AOI22_X1 p7_mult_21_U454 ( .A1(reg2_reg[11]), .A2(p7_mult_21_n885), .B1(
        B1[12]), .B2(p7_mult_21_n911), .ZN(p7_mult_21_n908) );
  AOI222_X1 p7_mult_21_U455 ( .A1(p7_mult_21_n916), .A2(p7_mult_21_n917), .B1(
        p7_mult_21_n916), .B2(p7_mult_21_n907), .C1(p7_mult_21_n917), .C2(
        p7_mult_21_n907), .ZN(p7_mult_21_n898) );
  OAI21_X1 p7_mult_21_U456 ( .B1(p7_mult_21_n919), .B2(p7_mult_21_n920), .A(
        p7_mult_21_n921), .ZN(p7_mult_21_n905) );
  AOI22_X1 p7_mult_21_U458 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n903), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n923), .ZN(p7_mult_21_n922) );
  OAI22_X1 p7_mult_21_U459 ( .A1(p7_mult_21_n876), .A2(B1[10]), .B1(
        p7_mult_21_n924), .B2(reg2_reg[13]), .ZN(p7_mult_21_n903) );
  XNOR2_X1 p7_mult_21_U466 ( .A(p7_mult_21_n938), .B(p7_mult_21_n930), .ZN(
        p7_mult_21_n927) );
  XNOR2_X1 p7_mult_21_U475 ( .A(p7_mult_21_n928), .B(p7_mult_21_n929), .ZN(
        p7_mult_21_n938) );
  AOI222_X1 p7_mult_21_U491 ( .A1(p7_mult_21_n975), .A2(p7_mult_21_n976), .B1(
        p7_mult_21_n975), .B2(p7_mult_21_n977), .C1(p7_mult_21_n976), .C2(
        p7_mult_21_n977), .ZN(p7_mult_21_n932) );
  XNOR2_X1 p7_mult_21_U495 ( .A(p7_mult_21_n985), .B(p7_mult_21_n977), .ZN(
        p7_mult_21_n974) );
  XNOR2_X1 p7_mult_21_U504 ( .A(p7_mult_21_n975), .B(p7_mult_21_n976), .ZN(
        p7_mult_21_n985) );
  XNOR2_X1 p7_mult_21_U505 ( .A(p7_mult_21_n963), .B(p7_mult_21_n995), .ZN(
        p7_mult_21_n976) );
  XNOR2_X1 p7_mult_21_U506 ( .A(p7_mult_21_n964), .B(p7_mult_21_n965), .ZN(
        p7_mult_21_n995) );
  AOI222_X1 p7_mult_21_U513 ( .A1(p7_mult_21_n1005), .A2(p7_mult_21_n1006), 
        .B1(p7_mult_21_n1005), .B2(p7_mult_21_n1007), .C1(p7_mult_21_n1006), 
        .C2(p7_mult_21_n1007), .ZN(p7_mult_21_n975) );
  AOI222_X1 p7_mult_21_U494 ( .A1(p7_mult_21_n982), .A2(p7_mult_21_n983), .B1(
        p7_mult_21_n982), .B2(p7_mult_21_n984), .C1(p7_mult_21_n983), .C2(
        p7_mult_21_n984), .ZN(p7_mult_21_n972) );
  AOI222_X1 p7_mult_21_U516 ( .A1(p7_mult_21_n1011), .A2(p7_mult_21_n1012), 
        .B1(p7_mult_21_n1011), .B2(p7_mult_21_n1013), .C1(p7_mult_21_n1012), 
        .C2(p7_mult_21_n1013), .ZN(p7_mult_21_n983) );
  AOI222_X1 p7_mult_21_U517 ( .A1(p7_mult_21_n1014), .A2(p7_mult_21_n1015), 
        .B1(p7_mult_21_n1014), .B2(p7_mult_21_n1016), .C1(p7_mult_21_n1015), 
        .C2(p7_mult_21_n1016), .ZN(p7_mult_21_n982) );
  XNOR2_X1 p7_mult_21_U518 ( .A(p7_mult_21_n1008), .B(p7_mult_21_n1006), .ZN(
        p7_mult_21_n1017) );
  OAI222_X1 p7_mult_21_U526 ( .A1(p7_mult_21_n1024), .A2(p7_mult_21_n1025), 
        .B1(p7_mult_21_n1024), .B2(p7_mult_21_n1026), .C1(p7_mult_21_n1025), 
        .C2(p7_mult_21_n1026), .ZN(p7_mult_21_n1008) );
  XNOR2_X1 p7_mult_21_U536 ( .A(p7_mult_21_n1047), .B(p7_mult_21_n1013), .ZN(
        p7_mult_21_n1038) );
  XNOR2_X1 p7_mult_21_U537 ( .A(p7_mult_21_n1025), .B(p7_mult_21_n1048), .ZN(
        p7_mult_21_n1013) );
  OAI22_X1 p7_mult_21_U538 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1023), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1049), .ZN(p7_mult_21_n1024) );
  OAI22_X1 p7_mult_21_U544 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n1019), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n1054), .ZN(p7_mult_21_n1025) );
  XNOR2_X1 p7_mult_21_U546 ( .A(p7_mult_21_n1011), .B(p7_mult_21_n1012), .ZN(
        p7_mult_21_n1047) );
  AOI222_X1 p7_mult_21_U547 ( .A1(p7_mult_21_n1055), .A2(p7_mult_21_n1056), 
        .B1(p7_mult_21_n1055), .B2(p7_mult_21_n1057), .C1(p7_mult_21_n1056), 
        .C2(p7_mult_21_n1057), .ZN(p7_mult_21_n1012) );
  AOI222_X1 p7_mult_21_U548 ( .A1(p7_mult_21_n1058), .A2(p7_mult_21_n1059), 
        .B1(p7_mult_21_n1058), .B2(p7_mult_21_n1060), .C1(p7_mult_21_n1059), 
        .C2(p7_mult_21_n1060), .ZN(p7_mult_21_n1011) );
  AOI222_X1 p7_mult_21_U550 ( .A1(p7_mult_21_n1062), .A2(p7_mult_21_n1063), 
        .B1(p7_mult_21_n1062), .B2(p7_mult_21_n1064), .C1(p7_mult_21_n1063), 
        .C2(p7_mult_21_n1064), .ZN(p7_mult_21_n1036) );
  XNOR2_X1 p7_mult_21_U551 ( .A(p7_mult_21_n1065), .B(p7_mult_21_n1016), .ZN(
        p7_mult_21_n1037) );
  AOI22_X1 p7_mult_21_U552 ( .A1(p7_mult_21_n919), .A2(p7_mult_21_n1021), .B1(
        p7_mult_21_n920), .B2(p7_mult_21_n1066), .ZN(p7_mult_21_n1016) );
  XNOR2_X1 p7_mult_21_U554 ( .A(p7_mult_21_n1014), .B(p7_mult_21_n1015), .ZN(
        p7_mult_21_n1065) );
  AOI22_X1 p7_mult_21_U555 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n1031), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n1067), .ZN(p7_mult_21_n1015) );
  AOI222_X1 p7_mult_21_U558 ( .A1(p7_mult_21_n1069), .A2(p7_mult_21_n1070), 
        .B1(p7_mult_21_n1069), .B2(p7_mult_21_n1071), .C1(p7_mult_21_n1070), 
        .C2(p7_mult_21_n1071), .ZN(p7_mult_21_n1014) );
  XNOR2_X1 p7_mult_21_U603 ( .A(p7_mult_21_n1104), .B(p7_mult_21_n1105), .ZN(
        p7_mult_21_n1114) );
  XNOR2_X1 p7_mult_21_U614 ( .A(p7_mult_21_n1119), .B(p7_mult_21_n1118), .ZN(
        p7_mult_21_n1154) );
  AOI222_X1 p7_mult_21_U622 ( .A1(p7_mult_21_n1163), .A2(p7_mult_21_n1164), 
        .B1(p7_mult_21_n1163), .B2(p7_mult_21_n1165), .C1(p7_mult_21_n1164), 
        .C2(p7_mult_21_n1165), .ZN(p7_mult_21_n1113) );
  XNOR2_X1 p7_mult_21_U623 ( .A(p7_mult_21_n1166), .B(p7_mult_21_n1145), .ZN(
        p7_mult_21_n1111) );
  XNOR2_X1 p7_mult_21_U630 ( .A(p7_mult_21_n1143), .B(p7_mult_21_n1144), .ZN(
        p7_mult_21_n1166) );
  AOI222_X1 p7_mult_21_U613 ( .A1(p7_mult_21_n1150), .A2(p7_mult_21_n1151), 
        .B1(p7_mult_21_n1150), .B2(p7_mult_21_n1152), .C1(p7_mult_21_n1151), 
        .C2(p7_mult_21_n1152), .ZN(p7_mult_21_n1110) );
  AOI222_X1 p7_mult_21_U755 ( .A1(p7_mult_21_n1188), .A2(p7_mult_21_n1189), 
        .B1(p7_mult_21_n1188), .B2(p7_mult_21_n1187), .C1(p7_mult_21_n1189), 
        .C2(p7_mult_21_n1187), .ZN(p7_mult_21_n1148) );
  XNOR2_X1 p7_mult_21_U777 ( .A(p7_mult_21_n1366), .B(p7_mult_21_n1163), .ZN(
        p7_mult_21_n1151) );
  AOI222_X1 p7_mult_21_U778 ( .A1(p7_mult_21_n1364), .A2(p7_mult_21_n1363), 
        .B1(p7_mult_21_n1364), .B2(p7_mult_21_n1367), .C1(p7_mult_21_n1363), 
        .C2(p7_mult_21_n1367), .ZN(p7_mult_21_n1163) );
  XNOR2_X1 p7_mult_21_U792 ( .A(p7_mult_21_n1164), .B(p7_mult_21_n1165), .ZN(
        p7_mult_21_n1366) );
  XNOR2_X1 p7_mult_21_U793 ( .A(p7_mult_21_n1375), .B(p7_mult_21_n1162), .ZN(
        p7_mult_21_n1165) );
  XNOR2_X1 p7_mult_21_U797 ( .A(p7_mult_21_n1160), .B(p7_mult_21_n1161), .ZN(
        p7_mult_21_n1375) );
  XNOR2_X1 p7_mult_21_U806 ( .A(p7_mult_21_n1159), .B(p7_mult_21_n1380), .ZN(
        p7_mult_21_n1164) );
  XNOR2_X1 p7_mult_21_U818 ( .A(p7_mult_21_n1384), .B(p7_mult_21_n1175), .ZN(
        p7_mult_21_n1152) );
  XNOR2_X1 p7_mult_21_U827 ( .A(p7_mult_21_n1174), .B(p7_mult_21_n1173), .ZN(
        p7_mult_21_n1384) );
  AOI222_X1 p7_mult_21_U830 ( .A1(p7_mult_21_n1358), .A2(p7_mult_21_n1360), 
        .B1(p7_mult_21_n1358), .B2(p7_mult_21_n1359), .C1(p7_mult_21_n1360), 
        .C2(p7_mult_21_n1359), .ZN(p7_mult_21_n1150) );
  XNOR2_X1 p7_mult_21_U639 ( .A(p7_mult_21_n1186), .B(p7_mult_21_n1187), .ZN(
        p7_mult_21_n1185) );
  AOI222_X1 p7_mult_21_U756 ( .A1(p7_mult_21_n1202), .A2(p7_mult_21_n1203), 
        .B1(p7_mult_21_n1202), .B2(p7_mult_21_n1201), .C1(p7_mult_21_n1203), 
        .C2(p7_mult_21_n1201), .ZN(p7_mult_21_n1187) );
  XNOR2_X1 p7_mult_21_U640 ( .A(p7_mult_21_n1188), .B(p7_mult_21_n1189), .ZN(
        p7_mult_21_n1186) );
  XNOR2_X1 p7_mult_21_U774 ( .A(p7_mult_21_n1357), .B(p7_mult_21_n1358), .ZN(
        p7_mult_21_n1189) );
  XNOR2_X1 p7_mult_21_U775 ( .A(p7_mult_21_n1359), .B(p7_mult_21_n1360), .ZN(
        p7_mult_21_n1357) );
  XNOR2_X1 p7_mult_21_U844 ( .A(p7_mult_21_n1399), .B(p7_mult_21_n1392), .ZN(
        p7_mult_21_n1360) );
  XNOR2_X1 p7_mult_21_U856 ( .A(p7_mult_21_n1390), .B(p7_mult_21_n1391), .ZN(
        p7_mult_21_n1399) );
  OAI222_X1 p7_mult_21_U831 ( .A1(p7_mult_21_n1205), .A2(p7_mult_21_n1207), 
        .B1(p7_mult_21_n1205), .B2(p7_mult_21_n1206), .C1(p7_mult_21_n1207), 
        .C2(p7_mult_21_n1206), .ZN(p7_mult_21_n1359) );
  XNOR2_X1 p7_mult_21_U776 ( .A(p7_mult_21_n1361), .B(p7_mult_21_n1362), .ZN(
        p7_mult_21_n1188) );
  NOR2_X1 p7_mult_21_U791 ( .A1(p7_mult_21_n1373), .A2(p7_mult_21_n1374), .ZN(
        p7_mult_21_n1364) );
  AOI222_X1 p7_mult_21_U781 ( .A1(p7_mult_21_n1347), .A2(p7_mult_21_n1348), 
        .B1(p7_mult_21_n1347), .B2(p7_mult_21_n1346), .C1(p7_mult_21_n1348), 
        .C2(p7_mult_21_n1346), .ZN(p7_mult_21_n1363) );
  AOI222_X1 p7_mult_21_U641 ( .A1(p7_mult_21_n1190), .A2(p7_mult_21_n1191), 
        .B1(p7_mult_21_n1190), .B2(p7_mult_21_n1192), .C1(p7_mult_21_n1191), 
        .C2(p7_mult_21_n1192), .ZN(p7_mult_21_n1184) );
  AOI222_X1 p7_mult_21_U643 ( .A1(p7_mult_21_n1196), .A2(p7_mult_21_n1197), 
        .B1(p7_mult_21_n1196), .B2(p7_mult_21_n1198), .C1(p7_mult_21_n1197), 
        .C2(p7_mult_21_n1198), .ZN(p7_mult_21_n1195) );
  XNOR2_X1 p7_mult_21_U644 ( .A(p7_mult_21_n1200), .B(p7_mult_21_n1201), .ZN(
        p7_mult_21_n1191) );
  XNOR2_X1 p7_mult_21_U757 ( .A(p7_mult_21_n1345), .B(p7_mult_21_n1346), .ZN(
        p7_mult_21_n1201) );
  AOI22_X1 p7_mult_21_U782 ( .A1(reg2_reg[0]), .A2(p7_mult_21_n1370), .B1(
        p7_mult_21_n1289), .B2(p7_mult_21_n1350), .ZN(p7_mult_21_n1346) );
  XNOR2_X1 p7_mult_21_U758 ( .A(p7_mult_21_n1347), .B(p7_mult_21_n1348), .ZN(
        p7_mult_21_n1345) );
  AOI22_X1 p7_mult_21_U787 ( .A1(reg2_reg[5]), .A2(B1[7]), .B1(p7_mult_21_n988), .B2(p7_mult_21_n1053), .ZN(p7_mult_21_n1369) );
  AOI22_X1 p7_mult_21_U788 ( .A1(p7_mult_21_n919), .A2(p7_mult_21_n1371), .B1(
        p7_mult_21_n920), .B2(p7_mult_21_n1356), .ZN(p7_mult_21_n1347) );
  XNOR2_X1 p7_mult_21_U645 ( .A(p7_mult_21_n1202), .B(p7_mult_21_n1203), .ZN(
        p7_mult_21_n1200) );
  AOI222_X1 p7_mult_21_U759 ( .A1(p7_mult_21_n1317), .A2(p7_mult_21_n1316), 
        .B1(p7_mult_21_n1317), .B2(p7_mult_21_n1315), .C1(p7_mult_21_n1316), 
        .C2(p7_mult_21_n1315), .ZN(p7_mult_21_n1203) );
  OAI222_X1 p7_mult_21_U766 ( .A1(p7_mult_21_n1323), .A2(p7_mult_21_n1324), 
        .B1(p7_mult_21_n1323), .B2(p7_mult_21_n1322), .C1(p7_mult_21_n1324), 
        .C2(p7_mult_21_n1322), .ZN(p7_mult_21_n1352) );
  XNOR2_X1 p7_mult_21_U646 ( .A(p7_mult_21_n1204), .B(p7_mult_21_n1205), .ZN(
        p7_mult_21_n1192) );
  XNOR2_X1 p7_mult_21_U839 ( .A(p7_mult_21_n1374), .B(p7_mult_21_n1373), .ZN(
        p7_mult_21_n1205) );
  AOI21_X1 p7_mult_21_U841 ( .B1(p7_mult_21_n1397), .B2(p7_mult_21_n886), .A(
        p7_mult_21_n1398), .ZN(p7_mult_21_n1374) );
  XNOR2_X1 p7_mult_21_U647 ( .A(p7_mult_21_n1206), .B(p7_mult_21_n1207), .ZN(
        p7_mult_21_n1204) );
  OAI22_X1 p7_mult_21_U833 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1394), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1351), .ZN(p7_mult_21_n1393) );
  AOI222_X1 p7_mult_21_U648 ( .A1(p7_mult_21_n1208), .A2(p7_mult_21_n1209), 
        .B1(p7_mult_21_n1208), .B2(p7_mult_21_n1210), .C1(p7_mult_21_n1209), 
        .C2(p7_mult_21_n1210), .ZN(p7_mult_21_n1190) );
  AOI222_X1 p7_mult_21_U652 ( .A1(p7_mult_21_n1218), .A2(p7_mult_21_n1219), 
        .B1(p7_mult_21_n1218), .B2(p7_mult_21_n1220), .C1(p7_mult_21_n1219), 
        .C2(p7_mult_21_n1220), .ZN(p7_mult_21_n1217) );
  XNOR2_X1 p7_mult_21_U654 ( .A(p7_mult_21_n1222), .B(p7_mult_21_n1223), .ZN(
        p7_mult_21_n1216) );
  XNOR2_X1 p7_mult_21_U655 ( .A(p7_mult_21_n1224), .B(p7_mult_21_n1225), .ZN(
        p7_mult_21_n1222) );
  XNOR2_X1 p7_mult_21_U697 ( .A(p7_mult_21_n1291), .B(p7_mult_21_n1292), .ZN(
        p7_mult_21_n1219) );
  XNOR2_X1 p7_mult_21_U698 ( .A(p7_mult_21_n1293), .B(p7_mult_21_n1294), .ZN(
        p7_mult_21_n1291) );
  AOI222_X1 p7_mult_21_U700 ( .A1(p7_mult_21_n1299), .A2(p7_mult_21_n1300), 
        .B1(p7_mult_21_n1299), .B2(p7_mult_21_n1301), .C1(p7_mult_21_n1300), 
        .C2(p7_mult_21_n1301), .ZN(p7_mult_21_n1221) );
  AOI222_X1 p7_mult_21_U701 ( .A1(p7_mult_21_n1237), .A2(p7_mult_21_n1235), 
        .B1(p7_mult_21_n1237), .B2(p7_mult_21_n1238), .C1(p7_mult_21_n1235), 
        .C2(p7_mult_21_n1238), .ZN(p7_mult_21_n1226) );
  XNOR2_X1 p7_mult_21_U702 ( .A(p7_mult_21_n1302), .B(p7_mult_21_n1303), .ZN(
        p7_mult_21_n1238) );
  XNOR2_X1 p7_mult_21_U703 ( .A(p7_mult_21_n1304), .B(p7_mult_21_n1301), .ZN(
        p7_mult_21_n1235) );
  OAI22_X1 p7_mult_21_U704 ( .A1(p7_mult_21_n1089), .A2(p7_mult_21_n1305), 
        .B1(p7_mult_21_n1051), .B2(p7_mult_21_n1279), .ZN(p7_mult_21_n1301) );
  AOI222_X1 p7_mult_21_U708 ( .A1(p7_mult_21_n1281), .A2(p7_mult_21_n1284), 
        .B1(p7_mult_21_n1281), .B2(p7_mult_21_n1283), .C1(p7_mult_21_n1284), 
        .C2(p7_mult_21_n1283), .ZN(p7_mult_21_n1237) );
  XNOR2_X1 p7_mult_21_U714 ( .A(p7_mult_21_n1310), .B(p7_mult_21_n1198), .ZN(
        p7_mult_21_n1213) );
  NOR2_X1 p7_mult_21_U715 ( .A1(p7_mult_21_n1312), .A2(p7_mult_21_n1313), .ZN(
        p7_mult_21_n1208) );
  XNOR2_X1 p7_mult_21_U716 ( .A(p7_mult_21_n1211), .B(p7_mult_21_n1209), .ZN(
        p7_mult_21_n1311) );
  XNOR2_X1 p7_mult_21_U717 ( .A(p7_mult_21_n1314), .B(p7_mult_21_n1315), .ZN(
        p7_mult_21_n1209) );
  NOR2_X1 p7_mult_21_U417 ( .A1(B1[9]), .A2(p7_mult_21_n1261), .ZN(
        p7_mult_21_n852) );
  XNOR2_X1 p7_mult_21_U718 ( .A(p7_mult_21_n1316), .B(p7_mult_21_n1317), .ZN(
        p7_mult_21_n1314) );
  OAI22_X1 p7_mult_21_U761 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1351), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1343), .ZN(p7_mult_21_n1316) );
  AOI222_X1 p7_mult_21_U719 ( .A1(p7_mult_21_n1318), .A2(p7_mult_21_n1319), 
        .B1(p7_mult_21_n1318), .B2(p7_mult_21_n1320), .C1(p7_mult_21_n1319), 
        .C2(p7_mult_21_n1320), .ZN(p7_mult_21_n1211) );
  XNOR2_X1 p7_mult_21_U720 ( .A(p7_mult_21_n1196), .B(p7_mult_21_n1197), .ZN(
        p7_mult_21_n1310) );
  XNOR2_X1 p7_mult_21_U721 ( .A(p7_mult_21_n1323), .B(p7_mult_21_n1324), .ZN(
        p7_mult_21_n1321) );
  AOI22_X1 p7_mult_21_U836 ( .A1(B1[8]), .A2(reg2_reg[3]), .B1(
        p7_mult_21_n1126), .B2(p7_mult_21_n962), .ZN(p7_mult_21_n1354) );
  AOI22_X1 p7_mult_21_U772 ( .A1(p7_mult_21_n919), .A2(p7_mult_21_n1356), .B1(
        n672), .B2(p7_mult_21_n1332), .ZN(p7_mult_21_n1323) );
  OAI222_X1 p7_mult_21_U722 ( .A1(p7_mult_21_n1325), .A2(p7_mult_21_n1326), 
        .B1(p7_mult_21_n1325), .B2(p7_mult_21_n1327), .C1(p7_mult_21_n1326), 
        .C2(p7_mult_21_n1327), .ZN(p7_mult_21_n1196) );
  AOI222_X1 p7_mult_21_U724 ( .A1(p7_mult_21_n1225), .A2(p7_mult_21_n1224), 
        .B1(p7_mult_21_n1225), .B2(p7_mult_21_n1223), .C1(p7_mult_21_n1224), 
        .C2(p7_mult_21_n1223), .ZN(p7_mult_21_n1212) );
  XNOR2_X1 p7_mult_21_U725 ( .A(p7_mult_21_n1329), .B(p7_mult_21_n1328), .ZN(
        p7_mult_21_n1223) );
  XNOR2_X1 p7_mult_21_U727 ( .A(p7_mult_21_n1313), .B(p7_mult_21_n1312), .ZN(
        p7_mult_21_n1325) );
  AOI21_X1 p7_mult_21_U729 ( .B1(p7_mult_21_n1332), .B2(p7_mult_21_n919), .A(
        p7_mult_21_n1333), .ZN(p7_mult_21_n1313) );
  AOI222_X1 p7_mult_21_U731 ( .A1(p7_mult_21_n1294), .A2(p7_mult_21_n1293), 
        .B1(p7_mult_21_n1294), .B2(p7_mult_21_n1292), .C1(p7_mult_21_n1293), 
        .C2(p7_mult_21_n1292), .ZN(p7_mult_21_n1327) );
  OAI22_X1 p7_mult_21_U733 ( .A1(p7_mult_21_n1089), .A2(p7_mult_21_n1335), 
        .B1(p7_mult_21_n1051), .B2(p7_mult_21_n1305), .ZN(p7_mult_21_n1293) );
  AOI222_X1 p7_mult_21_U736 ( .A1(p7_mult_21_n1298), .A2(p7_mult_21_n1297), 
        .B1(p7_mult_21_n1298), .B2(p7_mult_21_n1295), .C1(p7_mult_21_n1297), 
        .C2(p7_mult_21_n1295), .ZN(p7_mult_21_n1224) );
  AOI22_X1 p7_mult_21_U738 ( .A1(reg2_reg[3]), .A2(p7_mult_21_n1068), .B1(
        B1[5]), .B2(p7_mult_21_n1126), .ZN(p7_mult_21_n1307) );
  OAI22_X1 p7_mult_21_U739 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1337), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1338), .ZN(p7_mult_21_n1297) );
  OAI21_X1 p7_mult_21_U741 ( .B1(p7_mult_21_n1338), .B2(p7_mult_21_n1022), .A(
        p7_mult_21_n1339), .ZN(p7_mult_21_n1303) );
  OAI22_X1 p7_mult_21_U745 ( .A1(p7_mult_21_n1089), .A2(p7_mult_21_n1341), 
        .B1(p7_mult_21_n1051), .B2(p7_mult_21_n1335), .ZN(p7_mult_21_n1320) );
  AOI22_X1 p7_mult_21_U768 ( .A1(reg2_reg[5]), .A2(B1[5]), .B1(
        p7_mult_21_n1068), .B2(p7_mult_21_n1053), .ZN(p7_mult_21_n1342) );
  XNOR2_X1 p7_mult_21_U750 ( .A(p7_mult_21_n1318), .B(p7_mult_21_n1319), .ZN(
        p7_mult_21_n1340) );
  OAI22_X1 p7_mult_21_U751 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1343), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1337), .ZN(p7_mult_21_n1319) );
  OAI22_X1 p7_mult_21_U771 ( .A1(p7_mult_21_n988), .A2(p7_mult_21_n1126), .B1(
        reg2_reg[3]), .B2(B1[7]), .ZN(p7_mult_21_n1344) );
  XNOR2_X1 p7_mult_21_U604 ( .A(p7_mult_21_n1134), .B(p7_mult_21_n1103), .ZN(
        p7_mult_21_n1105) );
  XNOR2_X1 p7_mult_21_U606 ( .A(p7_mult_21_n1101), .B(p7_mult_21_n1102), .ZN(
        p7_mult_21_n1134) );
  AOI222_X1 p7_mult_21_U609 ( .A1(p7_mult_21_n1143), .A2(p7_mult_21_n1144), 
        .B1(p7_mult_21_n1143), .B2(p7_mult_21_n1145), .C1(p7_mult_21_n1144), 
        .C2(p7_mult_21_n1145), .ZN(p7_mult_21_n1104) );
  AOI222_X1 p7_mult_21_U631 ( .A1(p7_mult_21_n1173), .A2(p7_mult_21_n1174), 
        .B1(p7_mult_21_n1173), .B2(p7_mult_21_n1175), .C1(p7_mult_21_n1174), 
        .C2(p7_mult_21_n1175), .ZN(p7_mult_21_n1144) );
  XNOR2_X1 p7_mult_21_U819 ( .A(p7_mult_21_n1177), .B(p7_mult_21_n1178), .ZN(
        p7_mult_21_n1175) );
  AOI222_X1 p7_mult_21_U829 ( .A1(p7_mult_21_n1390), .A2(p7_mult_21_n1391), 
        .B1(p7_mult_21_n1390), .B2(p7_mult_21_n1392), .C1(p7_mult_21_n1391), 
        .C2(p7_mult_21_n1392), .ZN(p7_mult_21_n1174) );
  OAI22_X1 p7_mult_21_U845 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1382), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1394), .ZN(p7_mult_21_n1392) );
  AOI22_X1 p7_mult_21_U846 ( .A1(reg2_reg[7]), .A2(p7_mult_21_n1068), .B1(
        B1[5]), .B2(p7_mult_21_n992), .ZN(p7_mult_21_n1394) );
  AOI22_X1 p7_mult_21_U858 ( .A1(B1[9]), .A2(p7_mult_21_n1126), .B1(
        reg2_reg[3]), .B2(p7_mult_21_n941), .ZN(p7_mult_21_n1396) );
  AOI22_X1 p7_mult_21_U869 ( .A1(p7_mult_21_n886), .A2(p7_mult_21_n1379), .B1(
        p7_mult_21_n887), .B2(p7_mult_21_n1397), .ZN(p7_mult_21_n1402) );
  AOI222_X1 p7_mult_21_U828 ( .A1(p7_mult_21_n1387), .A2(p7_mult_21_n1388), 
        .B1(p7_mult_21_n1387), .B2(p7_mult_21_n1389), .C1(p7_mult_21_n1388), 
        .C2(p7_mult_21_n1389), .ZN(p7_mult_21_n1173) );
  OAI22_X1 p7_mult_21_U877 ( .A1(p7_mult_21_n970), .A2(p7_mult_21_n1377), .B1(
        p7_mult_21_n943), .B2(p7_mult_21_n1372), .ZN(p7_mult_21_n1388) );
  AOI222_X1 p7_mult_21_U535 ( .A1(p7_mult_21_n1043), .A2(p7_mult_21_n1044), 
        .B1(p7_mult_21_n1043), .B2(p7_mult_21_n1045), .C1(p7_mult_21_n1044), 
        .C2(p7_mult_21_n1045), .ZN(p7_mult_21_n1033) );
  OAI22_X1 p7_mult_21_U568 ( .A1(p7_mult_21_n1089), .A2(p7_mult_21_n1050), 
        .B1(p7_mult_21_n1051), .B2(p7_mult_21_n1090), .ZN(p7_mult_21_n1056) );
  OAI22_X1 p7_mult_21_U570 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n1054), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n1091), .ZN(p7_mult_21_n1055) );
  OAI22_X1 p7_mult_21_U572 ( .A1(p7_mult_21_n970), .A2(p7_mult_21_n1092), .B1(
        p7_mult_21_n943), .B2(p7_mult_21_n1093), .ZN(p7_mult_21_n1057) );
  AOI22_X1 p7_mult_21_U574 ( .A1(reg2_reg[9]), .A2(B1[8]), .B1(p7_mult_21_n962), .B2(p7_mult_21_n945), .ZN(p7_mult_21_n1066) );
  OAI22_X1 p7_mult_21_U576 ( .A1(p7_mult_21_n883), .A2(p7_mult_21_n1098), .B1(
        p7_mult_21_n874), .B2(p7_mult_21_n1099), .ZN(p7_mult_21_n1070) );
  AOI222_X1 p7_mult_21_U579 ( .A1(p7_mult_21_n1101), .A2(p7_mult_21_n1102), 
        .B1(p7_mult_21_n1101), .B2(p7_mult_21_n1103), .C1(p7_mult_21_n1102), 
        .C2(p7_mult_21_n1103), .ZN(p7_mult_21_n1062) );
  AOI222_X1 p7_mult_21_U607 ( .A1(p7_mult_21_n1137), .A2(p7_mult_21_n1138), 
        .B1(p7_mult_21_n1137), .B2(p7_mult_21_n1139), .C1(p7_mult_21_n1138), 
        .C2(p7_mult_21_n1139), .ZN(p7_mult_21_n1102) );
  OAI22_X1 p7_mult_21_U624 ( .A1(p7_mult_21_n970), .A2(p7_mult_21_n1130), .B1(
        p7_mult_21_n943), .B2(p7_mult_21_n1168), .ZN(p7_mult_21_n1138) );
  AOI222_X1 p7_mult_21_U608 ( .A1(p7_mult_21_n1140), .A2(p7_mult_21_n1141), 
        .B1(p7_mult_21_n1140), .B2(p7_mult_21_n1142), .C1(p7_mult_21_n1141), 
        .C2(p7_mult_21_n1142), .ZN(p7_mult_21_n1101) );
  OAI22_X1 p7_mult_21_U635 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1131), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1181), .ZN(p7_mult_21_n1142) );
  OAI22_X1 p7_mult_21_U633 ( .A1(p7_mult_21_n883), .A2(p7_mult_21_n1132), .B1(
        p7_mult_21_n874), .B2(p7_mult_21_n1179), .ZN(p7_mult_21_n1141) );
  OAI21_X1 p7_mult_21_U820 ( .B1(p7_mult_21_n1179), .B2(p7_mult_21_n883), .A(
        p7_mult_21_n1385), .ZN(p7_mult_21_n1178) );
  XNOR2_X1 p7_mult_21_U562 ( .A(p7_mult_21_n1058), .B(p7_mult_21_n1061), .ZN(
        p7_mult_21_n1077) );
  OAI222_X1 p7_mult_21_U563 ( .A1(p7_mult_21_n1078), .A2(p7_mult_21_n1079), 
        .B1(p7_mult_21_n1078), .B2(p7_mult_21_n1080), .C1(p7_mult_21_n1079), 
        .C2(p7_mult_21_n1080), .ZN(p7_mult_21_n1061) );
  AOI222_X1 p7_mult_21_U564 ( .A1(p7_mult_21_n1081), .A2(p7_mult_21_n1082), 
        .B1(p7_mult_21_n1081), .B2(p7_mult_21_n1071), .C1(p7_mult_21_n1082), 
        .C2(p7_mult_21_n1071), .ZN(p7_mult_21_n1058) );
  OAI22_X1 p7_mult_21_U565 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1049), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1083), .ZN(p7_mult_21_n1060) );
  OAI22_X1 p7_mult_21_U566 ( .A1(p7_mult_21_n992), .A2(p7_mult_21_n924), .B1(
        B1[10]), .B2(reg2_reg[7]), .ZN(p7_mult_21_n1049) );
  AOI222_X1 p7_mult_21_U567 ( .A1(p7_mult_21_n1084), .A2(p7_mult_21_n1085), 
        .B1(p7_mult_21_n1084), .B2(p7_mult_21_n1086), .C1(p7_mult_21_n1085), 
        .C2(p7_mult_21_n1086), .ZN(p7_mult_21_n1043) );
  OAI22_X1 p7_mult_21_U596 ( .A1(p7_mult_21_n970), .A2(p7_mult_21_n1093), .B1(
        p7_mult_21_n943), .B2(p7_mult_21_n1130), .ZN(p7_mult_21_n1080) );
  OAI22_X1 p7_mult_21_U597 ( .A1(p7_mult_21_n945), .A2(p7_mult_21_n988), .B1(
        B1[7]), .B2(reg2_reg[9]), .ZN(p7_mult_21_n1093) );
  XNOR2_X1 p7_mult_21_U598 ( .A(p7_mult_21_n1078), .B(p7_mult_21_n1079), .ZN(
        p7_mult_21_n1129) );
  OAI22_X1 p7_mult_21_U599 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1083), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1131), .ZN(p7_mult_21_n1079) );
  OAI22_X1 p7_mult_21_U636 ( .A1(p7_mult_21_n992), .A2(p7_mult_21_n962), .B1(
        B1[8]), .B2(reg2_reg[7]), .ZN(p7_mult_21_n1131) );
  OAI22_X1 p7_mult_21_U600 ( .A1(p7_mult_21_n992), .A2(p7_mult_21_n941), .B1(
        B1[9]), .B2(reg2_reg[7]), .ZN(p7_mult_21_n1083) );
  OAI22_X1 p7_mult_21_U601 ( .A1(p7_mult_21_n883), .A2(p7_mult_21_n1099), .B1(
        p7_mult_21_n874), .B2(p7_mult_21_n1132), .ZN(p7_mult_21_n1078) );
  OAI22_X1 p7_mult_21_U589 ( .A1(p7_mult_21_n904), .A2(p7_mult_21_n1053), .B1(
        reg2_reg[5]), .B2(B1[11]), .ZN(p7_mult_21_n1090) );
  AOI22_X1 p7_mult_21_U592 ( .A1(B1[13]), .A2(reg2_reg[3]), .B1(
        p7_mult_21_n1126), .B2(p7_mult_21_n877), .ZN(p7_mult_21_n1097) );
  AOI22_X1 p7_mult_21_U627 ( .A1(B1[12]), .A2(p7_mult_21_n1126), .B1(
        reg2_reg[3]), .B2(p7_mult_21_n885), .ZN(p7_mult_21_n1123) );
  AOI22_X1 p7_mult_21_U593 ( .A1(p7_mult_21_n886), .A2(p7_mult_21_n1127), .B1(
        n673), .B2(p7_mult_21_n1128), .ZN(p7_mult_21_n1082) );
  OAI22_X1 p7_mult_21_U595 ( .A1(p7_mult_21_n911), .A2(p7_mult_21_n1068), .B1(
        B1[5]), .B2(reg2_reg[11]), .ZN(p7_mult_21_n1091) );
  AOI222_X1 p7_mult_21_U585 ( .A1(p7_mult_21_n1116), .A2(p7_mult_21_n1117), 
        .B1(p7_mult_21_n1116), .B2(p7_mult_21_n1118), .C1(p7_mult_21_n1117), 
        .C2(p7_mult_21_n1118), .ZN(p7_mult_21_n1084) );
  XNOR2_X1 p7_mult_21_U615 ( .A(p7_mult_21_n1135), .B(p7_mult_21_n1136), .ZN(
        p7_mult_21_n1118) );
  AOI22_X1 p7_mult_21_U616 ( .A1(p7_mult_21_n886), .A2(p7_mult_21_n1128), .B1(
        p7_mult_21_n887), .B2(p7_mult_21_n1155), .ZN(p7_mult_21_n1136) );
  AOI22_X1 p7_mult_21_U619 ( .A1(B1[10]), .A2(reg2_reg[5]), .B1(
        p7_mult_21_n1053), .B2(p7_mult_21_n924), .ZN(p7_mult_21_n1122) );
  AOI222_X1 p7_mult_21_U621 ( .A1(p7_mult_21_n1160), .A2(p7_mult_21_n1161), 
        .B1(p7_mult_21_n1160), .B2(p7_mult_21_n1162), .C1(p7_mult_21_n1161), 
        .C2(p7_mult_21_n1162), .ZN(p7_mult_21_n1117) );
  OAI22_X1 p7_mult_21_U795 ( .A1(p7_mult_21_n970), .A2(p7_mult_21_n1168), .B1(
        p7_mult_21_n943), .B2(p7_mult_21_n1377), .ZN(p7_mult_21_n1376) );
  AOI22_X1 p7_mult_21_U796 ( .A1(reg2_reg[9]), .A2(p7_mult_21_n1068), .B1(
        B1[5]), .B2(p7_mult_21_n945), .ZN(p7_mult_21_n1168) );
  AOI22_X1 p7_mult_21_U799 ( .A1(B1[8]), .A2(reg2_reg[5]), .B1(
        p7_mult_21_n1053), .B2(p7_mult_21_n962), .ZN(p7_mult_21_n1368) );
  OAI22_X1 p7_mult_21_U801 ( .A1(p7_mult_21_n941), .A2(reg2_reg[5]), .B1(
        p7_mult_21_n1053), .B2(B1[9]), .ZN(p7_mult_21_n1156) );
  AOI22_X1 p7_mult_21_U804 ( .A1(p7_mult_21_n886), .A2(p7_mult_21_n1155), .B1(
        p7_mult_21_n887), .B2(p7_mult_21_n1379), .ZN(p7_mult_21_n1160) );
  OAI222_X1 p7_mult_21_U620 ( .A1(p7_mult_21_n1157), .A2(p7_mult_21_n1158), 
        .B1(p7_mult_21_n1157), .B2(p7_mult_21_n1159), .C1(p7_mult_21_n1158), 
        .C2(p7_mult_21_n1159), .ZN(p7_mult_21_n1119) );
  OAI22_X1 p7_mult_21_U862 ( .A1(p7_mult_21_n924), .A2(p7_mult_21_n1126), .B1(
        reg2_reg[3]), .B2(B1[10]), .ZN(p7_mult_21_n1383) );
  AOI22_X1 p7_mult_21_U816 ( .A1(B1[11]), .A2(p7_mult_21_n1126), .B1(
        reg2_reg[3]), .B2(p7_mult_21_n904), .ZN(p7_mult_21_n1170) );
  OAI22_X1 p7_mult_21_U812 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n1181), 
        .B1(p7_mult_21_n990), .B2(p7_mult_21_n1382), .ZN(p7_mult_21_n1158) );
  AOI22_X1 p7_mult_21_U813 ( .A1(reg2_reg[7]), .A2(p7_mult_21_n988), .B1(B1[7]), .B2(p7_mult_21_n992), .ZN(p7_mult_21_n1181) );
  OAI22_X1 p7_mult_21_U807 ( .A1(p7_mult_21_n1260), .A2(p7_mult_21_n1172), 
        .B1(p7_mult_21_n1271), .B2(p7_mult_21_n1381), .ZN(p7_mult_21_n1157) );
  NOR2_X1 p7_mult_21_U809 ( .A1(reg2_reg[0]), .A2(p7_mult_21_n1261), .ZN(
        p7_mult_21_n1289) );
  AOI222_X1 p7_mult_21_U465 ( .A1(p7_mult_21_n935), .A2(p7_mult_21_n936), .B1(
        p7_mult_21_n935), .B2(p7_mult_21_n937), .C1(p7_mult_21_n936), .C2(
        p7_mult_21_n937), .ZN(p7_mult_21_n925) );
  AOI222_X1 p7_mult_21_U483 ( .A1(p7_mult_21_n963), .A2(p7_mult_21_n964), .B1(
        p7_mult_21_n963), .B2(p7_mult_21_n965), .C1(p7_mult_21_n964), .C2(
        p7_mult_21_n965), .ZN(p7_mult_21_n935) );
  AOI22_X1 p7_mult_21_U507 ( .A1(p7_mult_21_n919), .A2(p7_mult_21_n996), .B1(
        p7_mult_21_n920), .B2(p7_mult_21_n997), .ZN(p7_mult_21_n965) );
  AOI222_X1 p7_mult_21_U510 ( .A1(p7_mult_21_n998), .A2(p7_mult_21_n999), .B1(
        p7_mult_21_n998), .B2(p7_mult_21_n1000), .C1(p7_mult_21_n999), .C2(
        p7_mult_21_n1000), .ZN(p7_mult_21_n964) );
  OAI21_X1 p7_mult_21_U541 ( .B1(p7_mult_21_n1050), .B2(p7_mult_21_n1051), .A(
        p7_mult_21_n1052), .ZN(p7_mult_21_n1000) );
  AOI22_X1 p7_mult_21_U569 ( .A1(B1[12]), .A2(p7_mult_21_n1053), .B1(
        reg2_reg[5]), .B2(p7_mult_21_n885), .ZN(p7_mult_21_n1050) );
  AOI22_X1 p7_mult_21_U528 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n987), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n1031), .ZN(p7_mult_21_n1001) );
  OAI22_X1 p7_mult_21_U556 ( .A1(p7_mult_21_n876), .A2(B1[5]), .B1(
        p7_mult_21_n1068), .B2(reg2_reg[13]), .ZN(p7_mult_21_n1031) );
  AOI22_X1 p7_mult_21_U543 ( .A1(B1[13]), .A2(reg2_reg[5]), .B1(
        p7_mult_21_n1053), .B2(p7_mult_21_n877), .ZN(p7_mult_21_n1030) );
  AOI222_X1 p7_mult_21_U512 ( .A1(p7_mult_21_n1002), .A2(p7_mult_21_n1003), 
        .B1(p7_mult_21_n1002), .B2(p7_mult_21_n1004), .C1(p7_mult_21_n1003), 
        .C2(p7_mult_21_n1004), .ZN(p7_mult_21_n963) );
  OAI22_X1 p7_mult_21_U524 ( .A1(p7_mult_21_n1022), .A2(p7_mult_21_n989), .B1(
        p7_mult_21_n990), .B2(p7_mult_21_n1023), .ZN(p7_mult_21_n1004) );
  AOI22_X1 p7_mult_21_U539 ( .A1(B1[11]), .A2(p7_mult_21_n992), .B1(
        reg2_reg[7]), .B2(p7_mult_21_n904), .ZN(p7_mult_21_n1023) );
  OAI22_X1 p7_mult_21_U519 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n994), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n1019), .ZN(p7_mult_21_n1003) );
  AOI22_X1 p7_mult_21_U545 ( .A1(reg2_reg[11]), .A2(p7_mult_21_n988), .B1(
        B1[7]), .B2(p7_mult_21_n911), .ZN(p7_mult_21_n1019) );
  AOI22_X1 p7_mult_21_U522 ( .A1(p7_mult_21_n919), .A2(p7_mult_21_n997), .B1(
        p7_mult_21_n920), .B2(p7_mult_21_n1021), .ZN(p7_mult_21_n1020) );
  OAI22_X1 p7_mult_21_U553 ( .A1(p7_mult_21_n945), .A2(B1[9]), .B1(
        p7_mult_21_n941), .B2(reg2_reg[9]), .ZN(p7_mult_21_n1021) );
  OAI22_X1 p7_mult_21_U523 ( .A1(p7_mult_21_n945), .A2(B1[10]), .B1(
        p7_mult_21_n924), .B2(reg2_reg[9]), .ZN(p7_mult_21_n997) );
  AOI22_X1 p7_mult_21_U467 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n923), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n940), .ZN(p7_mult_21_n916) );
  OAI22_X1 p7_mult_21_U468 ( .A1(p7_mult_21_n876), .A2(B1[9]), .B1(
        p7_mult_21_n941), .B2(reg2_reg[13]), .ZN(p7_mult_21_n923) );
  OAI21_X1 p7_mult_21_U469 ( .B1(p7_mult_21_n942), .B2(p7_mult_21_n943), .A(
        p7_mult_21_n944), .ZN(p7_mult_21_n907) );
  NAND2_X1 p7_mult_21_U470 ( .A1(p7_mult_21_n919), .A2(p7_mult_21_n921), .ZN(
        p7_mult_21_n944) );
  AOI22_X1 p7_mult_21_U471 ( .A1(B1[13]), .A2(reg2_reg[9]), .B1(
        p7_mult_21_n945), .B2(p7_mult_21_n877), .ZN(p7_mult_21_n921) );
  OAI22_X1 p7_mult_21_U473 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n915), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n947), .ZN(p7_mult_21_n946) );
  OAI22_X1 p7_mult_21_U474 ( .A1(p7_mult_21_n911), .A2(p7_mult_21_n904), .B1(
        B1[11]), .B2(reg2_reg[11]), .ZN(p7_mult_21_n915) );
  AOI222_X1 p7_mult_21_U476 ( .A1(p7_mult_21_n948), .A2(p7_mult_21_n949), .B1(
        p7_mult_21_n948), .B2(p7_mult_21_n950), .C1(p7_mult_21_n949), .C2(
        p7_mult_21_n950), .ZN(p7_mult_21_n929) );
  OAI22_X1 p7_mult_21_U487 ( .A1(p7_mult_21_n970), .A2(p7_mult_21_n942), .B1(
        p7_mult_21_n943), .B2(p7_mult_21_n971), .ZN(p7_mult_21_n950) );
  AOI22_X1 p7_mult_21_U509 ( .A1(reg2_reg[9]), .A2(p7_mult_21_n904), .B1(
        B1[11]), .B2(p7_mult_21_n945), .ZN(p7_mult_21_n971) );
  AOI22_X1 p7_mult_21_U488 ( .A1(B1[12]), .A2(p7_mult_21_n945), .B1(
        reg2_reg[9]), .B2(p7_mult_21_n885), .ZN(p7_mult_21_n942) );
  OAI22_X1 p7_mult_21_U484 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n947), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n967), .ZN(p7_mult_21_n949) );
  OAI22_X1 p7_mult_21_U485 ( .A1(p7_mult_21_n911), .A2(p7_mult_21_n924), .B1(
        B1[10]), .B2(reg2_reg[11]), .ZN(p7_mult_21_n947) );
  AOI222_X1 p7_mult_21_U486 ( .A1(p7_mult_21_n968), .A2(p7_mult_21_n969), .B1(
        p7_mult_21_n968), .B2(p7_mult_21_n953), .C1(p7_mult_21_n969), .C2(
        p7_mult_21_n953), .ZN(p7_mult_21_n948) );
  OAI22_X1 p7_mult_21_U502 ( .A1(p7_mult_21_n914), .A2(p7_mult_21_n967), .B1(
        p7_mult_21_n909), .B2(p7_mult_21_n994), .ZN(p7_mult_21_n993) );
  OAI22_X1 p7_mult_21_U520 ( .A1(p7_mult_21_n911), .A2(p7_mult_21_n962), .B1(
        B1[8]), .B2(reg2_reg[11]), .ZN(p7_mult_21_n994) );
  OAI22_X1 p7_mult_21_U503 ( .A1(p7_mult_21_n911), .A2(p7_mult_21_n941), .B1(
        B1[9]), .B2(reg2_reg[11]), .ZN(p7_mult_21_n967) );
  AOI22_X1 p7_mult_21_U496 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n961), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n987), .ZN(p7_mult_21_n968) );
  AOI222_X1 p7_mult_21_U477 ( .A1(p7_mult_21_n951), .A2(p7_mult_21_n952), .B1(
        p7_mult_21_n951), .B2(p7_mult_21_n953), .C1(p7_mult_21_n952), .C2(
        p7_mult_21_n953), .ZN(p7_mult_21_n928) );
  OAI21_X1 p7_mult_21_U498 ( .B1(p7_mult_21_n989), .B2(p7_mult_21_n990), .A(
        p7_mult_21_n991), .ZN(p7_mult_21_n953) );
  NAND2_X1 p7_mult_21_U499 ( .A1(p7_mult_21_n957), .A2(p7_mult_21_n959), .ZN(
        p7_mult_21_n991) );
  AOI22_X1 p7_mult_21_U525 ( .A1(B1[12]), .A2(p7_mult_21_n992), .B1(
        reg2_reg[7]), .B2(p7_mult_21_n885), .ZN(p7_mult_21_n989) );
  AOI22_X1 p7_mult_21_U481 ( .A1(p7_mult_21_n866), .A2(p7_mult_21_n940), .B1(
        p7_mult_21_n867), .B2(p7_mult_21_n961), .ZN(p7_mult_21_n960) );
  OAI22_X1 p7_mult_21_U497 ( .A1(p7_mult_21_n876), .A2(B1[7]), .B1(
        p7_mult_21_n988), .B2(reg2_reg[13]), .ZN(p7_mult_21_n961) );
  OAI221_X1 p7_mult_21_U825 ( .B1(reg2_reg[12]), .B2(reg2_reg[13]), .C1(
        p7_mult_21_n1386), .C2(p7_mult_21_n876), .A(p7_mult_21_n883), .ZN(
        p7_mult_21_n874) );
  AOI22_X1 p7_mult_21_U482 ( .A1(reg2_reg[13]), .A2(B1[8]), .B1(
        p7_mult_21_n962), .B2(p7_mult_21_n876), .ZN(p7_mult_21_n940) );
  OAI21_X1 p7_mult_21_U479 ( .B1(p7_mult_21_n957), .B2(p7_mult_21_n958), .A(
        p7_mult_21_n959), .ZN(p7_mult_21_n951) );
  AOI22_X1 p7_mult_21_U500 ( .A1(B1[13]), .A2(reg2_reg[7]), .B1(
        p7_mult_21_n992), .B2(p7_mult_21_n877), .ZN(p7_mult_21_n959) );
  AOI221_X1 p7_mult_21_U849 ( .B1(reg2_reg[6]), .B2(reg2_reg[7]), .C1(
        p7_mult_21_n1400), .C2(p7_mult_21_n992), .A(p7_mult_21_n957), .ZN(
        p7_mult_21_n958) );
  AOI22_X1 p7_mult_21_U853 ( .A1(reg2_reg[6]), .A2(reg2_reg[5]), .B1(
        p7_mult_21_n1053), .B2(p7_mult_21_n1400), .ZN(p7_mult_21_n957) );
  XOR2_X1 p7_mult_21_U983 ( .A(p7_mult_21_n1387), .B(p7_mult_21_n1388), .Z(
        p7_mult_21_n1404) );
  XOR2_X1 p7_mult_21_U982 ( .A(p7_mult_21_n1389), .B(p7_mult_21_n1404), .Z(
        p7_mult_21_n1358) );
  XOR2_X1 p7_mult_21_U981 ( .A(p7_mult_21_n1150), .B(p7_mult_21_n1152), .Z(
        p7_mult_21_n1365) );
  XOR2_X1 p7_mult_21_U980 ( .A(p7_mult_21_n1158), .B(p7_mult_21_n1157), .Z(
        p7_mult_21_n1380) );
  XOR2_X1 p7_mult_21_U979 ( .A(p7_mult_21_n1365), .B(p7_mult_21_n1151), .Z(
        p7_mult_21_n1149) );
  XOR2_X1 p7_mult_21_U978 ( .A(p7_mult_21_n1363), .B(p7_mult_21_n1364), .Z(
        p7_mult_21_n1362) );
  XOR2_X1 p7_mult_21_U977 ( .A(p7_mult_21_n1340), .B(p7_mult_21_n1320), .Z(
        p7_mult_21_n1225) );
  XOR2_X1 p7_mult_21_U976 ( .A(p7_mult_21_n1327), .B(p7_mult_21_n1325), .Z(
        p7_mult_21_n1329) );
  XOR2_X1 p7_mult_21_U975 ( .A(p7_mult_21_n1321), .B(p7_mult_21_n1322), .Z(
        p7_mult_21_n1197) );
  XOR2_X1 p7_mult_21_U974 ( .A(p7_mult_21_n1311), .B(p7_mult_21_n1208), .Z(
        p7_mult_21_n1198) );
  XOR2_X1 p7_mult_21_U973 ( .A(p7_mult_21_n1299), .B(p7_mult_21_n1300), .Z(
        p7_mult_21_n1304) );
  XOR2_X1 p7_mult_21_U972 ( .A(p7_mult_21_n1297), .B(p7_mult_21_n1298), .Z(
        p7_mult_21_n1296) );
  XOR2_X1 p7_mult_21_U971 ( .A(p7_mult_21_n1295), .B(p7_mult_21_n1296), .Z(
        p7_mult_21_n1218) );
  XOR2_X1 p7_mult_21_U970 ( .A(p7_mult_21_n1290), .B(p7_mult_21_n1219), .Z(
        p7_mult_21_n1227) );
  XOR2_X1 p7_mult_21_U965 ( .A(p7_mult_21_n1237), .B(p7_mult_21_n1238), .Z(
        p7_mult_21_n1236) );
  XOR2_X1 p7_mult_21_U964 ( .A(p7_mult_21_n1235), .B(p7_mult_21_n1236), .Z(
        p7_mult_21_n1230) );
  XOR2_X1 p7_mult_21_U963 ( .A(p7_mult_21_n1190), .B(p7_mult_21_n1192), .Z(
        p7_mult_21_n1199) );
  XOR2_X1 p7_mult_21_U962 ( .A(p7_mult_21_n1199), .B(p7_mult_21_n1191), .Z(
        p7_mult_21_n1194) );
  XOR2_X1 p7_mult_21_U961 ( .A(p7_mult_21_n1148), .B(p7_mult_21_n1147), .Z(
        p7_mult_21_n1182) );
  XOR2_X1 p7_mult_21_U960 ( .A(p7_mult_21_n1141), .B(p7_mult_21_n1140), .Z(
        p7_mult_21_n1176) );
  XOR2_X1 p7_mult_21_U959 ( .A(p7_mult_21_n1142), .B(p7_mult_21_n1176), .Z(
        p7_mult_21_n1143) );
  XOR2_X1 p7_mult_21_U958 ( .A(p7_mult_21_n1139), .B(p7_mult_21_n1138), .Z(
        p7_mult_21_n1167) );
  XOR2_X1 p7_mult_21_U957 ( .A(p7_mult_21_n1137), .B(p7_mult_21_n1167), .Z(
        p7_mult_21_n1145) );
  XOR2_X1 p7_mult_21_U956 ( .A(p7_mult_21_n1117), .B(p7_mult_21_n1154), .Z(
        p7_mult_21_n1112) );
  XOR2_X1 p7_mult_21_U955 ( .A(p7_mult_21_n1113), .B(p7_mult_21_n1112), .Z(
        p7_mult_21_n1153) );
  XOR2_X1 p7_mult_21_U954 ( .A(p7_mult_21_n1111), .B(p7_mult_21_n1153), .Z(
        p7_mult_21_n1108) );
  XOR2_X1 p7_mult_21_U953 ( .A(p7_mult_21_n1129), .B(p7_mult_21_n1080), .Z(
        p7_mult_21_n1086) );
  XOR2_X1 p7_mult_21_U952 ( .A(p7_mult_21_n1071), .B(p7_mult_21_n1081), .Z(
        p7_mult_21_n1120) );
  XOR2_X1 p7_mult_21_U951 ( .A(p7_mult_21_n1082), .B(p7_mult_21_n1120), .Z(
        p7_mult_21_n1085) );
  XOR2_X1 p7_mult_21_U950 ( .A(p7_mult_21_n1085), .B(p7_mult_21_n1084), .Z(
        p7_mult_21_n1115) );
  XOR2_X1 p7_mult_21_U949 ( .A(p7_mult_21_n1086), .B(p7_mult_21_n1115), .Z(
        p7_mult_21_n1106) );
  XOR2_X1 p7_mult_21_U948 ( .A(p7_mult_21_n1073), .B(p7_mult_21_n1074), .Z(
        p7_mult_21_n1107) );
  XOR2_X1 p7_mult_21_U947 ( .A(p7_mult_21_n1071), .B(p7_mult_21_n1070), .Z(
        p7_mult_21_n1094) );
  XOR2_X1 p7_mult_21_U946 ( .A(p7_mult_21_n1094), .B(p7_mult_21_n1069), .Z(
        p7_mult_21_n1063) );
  XOR2_X1 p7_mult_21_U945 ( .A(p7_mult_21_n1055), .B(p7_mult_21_n1056), .Z(
        p7_mult_21_n1088) );
  XOR2_X1 p7_mult_21_U944 ( .A(p7_mult_21_n1057), .B(p7_mult_21_n1088), .Z(
        p7_mult_21_n1064) );
  XOR2_X1 p7_mult_21_U943 ( .A(p7_mult_21_n1063), .B(p7_mult_21_n1064), .Z(
        p7_mult_21_n1087) );
  XOR2_X1 p7_mult_21_U942 ( .A(p7_mult_21_n1062), .B(p7_mult_21_n1087), .Z(
        p7_mult_21_n1045) );
  XOR2_X1 p7_mult_21_U941 ( .A(p7_mult_21_n1060), .B(p7_mult_21_n1077), .Z(
        p7_mult_21_n1044) );
  XOR2_X1 p7_mult_21_U940 ( .A(p7_mult_21_n1043), .B(p7_mult_21_n1044), .Z(
        p7_mult_21_n1076) );
  XOR2_X1 p7_mult_21_U939 ( .A(p7_mult_21_n1045), .B(p7_mult_21_n1076), .Z(
        p7_mult_21_n1041) );
  XOR2_X1 p7_mult_21_U938 ( .A(p7_mult_21_n1026), .B(p7_mult_21_n1024), .Z(
        p7_mult_21_n1048) );
  XOR2_X1 p7_mult_21_U937 ( .A(p7_mult_21_n1036), .B(p7_mult_21_n1038), .Z(
        p7_mult_21_n1046) );
  XOR2_X1 p7_mult_21_U936 ( .A(p7_mult_21_n1037), .B(p7_mult_21_n1046), .Z(
        p7_mult_21_n1035) );
  XOR2_X1 p7_mult_21_U935 ( .A(p7_mult_21_n1033), .B(n821), .Z(
        p7_mult_21_n1039) );
  XOR2_X1 p7_mult_21_U934 ( .A(p7_mult_21_n1026), .B(p7_mult_21_n1001), .Z(
        p7_mult_21_n1027) );
  XOR2_X1 p7_mult_21_U933 ( .A(p7_mult_21_n1027), .B(p7_mult_21_n998), .Z(
        p7_mult_21_n1007) );
  XOR2_X1 p7_mult_21_U932 ( .A(p7_mult_21_n1002), .B(p7_mult_21_n1003), .Z(
        p7_mult_21_n1018) );
  XOR2_X1 p7_mult_21_U931 ( .A(p7_mult_21_n1004), .B(p7_mult_21_n1018), .Z(
        p7_mult_21_n1006) );
  XOR2_X1 p7_mult_21_U930 ( .A(p7_mult_21_n1007), .B(p7_mult_21_n1017), .Z(
        p7_mult_21_n984) );
  XOR2_X1 p7_mult_21_U929 ( .A(p7_mult_21_n982), .B(p7_mult_21_n983), .Z(
        p7_mult_21_n1010) );
  XOR2_X1 p7_mult_21_U928 ( .A(p7_mult_21_n984), .B(p7_mult_21_n1010), .Z(
        p7_mult_21_n981) );
  XOR2_X1 p7_mult_21_U927 ( .A(p7_mult_21_n953), .B(p7_mult_21_n968), .Z(
        p7_mult_21_n986) );
  XOR2_X1 p7_mult_21_U926 ( .A(p7_mult_21_n969), .B(p7_mult_21_n986), .Z(
        p7_mult_21_n977) );
  XOR2_X1 p7_mult_21_U925 ( .A(p7_mult_21_n972), .B(n832), .Z(p7_mult_21_n978)
         );
  XOR2_X1 p7_mult_21_U924 ( .A(p7_mult_21_n948), .B(p7_mult_21_n949), .Z(
        p7_mult_21_n966) );
  XOR2_X1 p7_mult_21_U923 ( .A(p7_mult_21_n950), .B(p7_mult_21_n966), .Z(
        p7_mult_21_n937) );
  XOR2_X1 p7_mult_21_U922 ( .A(p7_mult_21_n953), .B(p7_mult_21_n952), .Z(
        p7_mult_21_n956) );
  XOR2_X1 p7_mult_21_U921 ( .A(p7_mult_21_n956), .B(p7_mult_21_n951), .Z(
        p7_mult_21_n936) );
  XOR2_X1 p7_mult_21_U920 ( .A(p7_mult_21_n935), .B(p7_mult_21_n936), .Z(
        p7_mult_21_n955) );
  XOR2_X1 p7_mult_21_U919 ( .A(p7_mult_21_n937), .B(p7_mult_21_n955), .Z(
        p7_mult_21_n934) );
  XOR2_X1 p7_mult_21_U918 ( .A(p7_mult_21_n907), .B(p7_mult_21_n916), .Z(
        p7_mult_21_n939) );
  XOR2_X1 p7_mult_21_U917 ( .A(p7_mult_21_n917), .B(p7_mult_21_n939), .Z(
        p7_mult_21_n930) );
  XOR2_X1 p7_mult_21_U916 ( .A(p7_mult_21_n925), .B(p7_mult_21_n926), .Z(
        p7_mult_21_n931) );
  XOR2_X1 p7_mult_21_U915 ( .A(p7_mult_21_n907), .B(p7_mult_21_n906), .Z(
        p7_mult_21_n918) );
  XOR2_X1 p7_mult_21_U914 ( .A(p7_mult_21_n918), .B(p7_mult_21_n905), .Z(
        p7_mult_21_n900) );
  XOR2_X1 p7_mult_21_U913 ( .A(p7_mult_21_n898), .B(p7_mult_21_n899), .Z(
        p7_mult_21_n913) );
  XOR2_X1 p7_mult_21_U911 ( .A(p7_mult_21_n872), .B(p7_mult_21_n892), .Z(
        p7_mult_21_n901) );
  XOR2_X1 p7_mult_21_U909 ( .A(p7_mult_21_n889), .B(n828), .Z(p7_mult_21_n894)
         );
  XOR2_X1 p7_mult_21_U908 ( .A(p7_mult_21_n872), .B(p7_mult_21_n871), .Z(
        p7_mult_21_n882) );
  XOR2_X1 p7_mult_21_U907 ( .A(p7_mult_21_n870), .B(p7_mult_21_n882), .Z(
        p7_mult_21_n880) );
  XOR2_X1 p7_mult_21_U906 ( .A(p7_mult_21_n860), .B(p7_mult_21_n864), .Z(
        p7_mult_21_n869) );
  MUX2_X1 p7_mult_21_U902 ( .A(p7_mult_21_n852), .B(p7_mult_21_n1350), .S(
        reg2_reg[0]), .Z(p7_mult_21_n1315) );
  INV_X1 p8_mult_21_U716 ( .A(p8_mult_21_n267), .ZN(p8_mult_21_n826) );
  INV_X1 p8_mult_21_U717 ( .A(p8_mult_21_n258), .ZN(p8_mult_21_n825) );
  INV_X1 p8_mult_21_U471 ( .A(p8_mult_21_n315), .ZN(p8_mult_21_n681) );
  INV_X1 p8_mult_21_U472 ( .A(p8_mult_21_n314), .ZN(p8_mult_21_n682) );
  INV_X1 p8_mult_21_U728 ( .A(B2[0]), .ZN(p8_mult_21_n721) );
  OR2_X1 p8_mult_21_U669 ( .A1(p8_mult_21_n816), .A2(p8_mult_21_n817), .ZN(
        p8_mult_21_n243) );
  INV_X1 p8_mult_21_U501 ( .A(p8_mult_21_n702), .ZN(p8_mult_21_n408) );
  INV_X1 p8_mult_21_U528 ( .A(p8_mult_21_n719), .ZN(p8_mult_21_n394) );
  INV_X1 p8_mult_21_U676 ( .A(p8_mult_21_n231), .ZN(p8_mult_21_n232) );
  INV_X1 p8_mult_21_U423 ( .A(p8_mult_21_n836), .ZN(p8_mult_21_n706) );
  INV_X1 p8_mult_21_U680 ( .A(p8_mult_21_n209), .ZN(p8_mult_21_n210) );
  INV_X1 p8_mult_21_U552 ( .A(p8_mult_21_n737), .ZN(p8_mult_21_n380) );
  NAND2_X1 p8_mult_21_U452 ( .A1(p8_mult_21_n722), .A2(p8_mult_21_n818), .ZN(
        p8_mult_21_n724) );
  INV_X1 p8_mult_21_U685 ( .A(p8_mult_21_n191), .ZN(p8_mult_21_n192) );
  INV_X1 p8_mult_21_U579 ( .A(p8_mult_21_n754), .ZN(p8_mult_21_n366) );
  NAND2_X1 p8_mult_21_U688 ( .A1(p8_mult_21_n739), .A2(p8_mult_21_n820), .ZN(
        p8_mult_21_n741) );
  INV_X1 p8_mult_21_U692 ( .A(p8_mult_21_n177), .ZN(p8_mult_21_n178) );
  INV_X1 p8_mult_21_U606 ( .A(p8_mult_21_n771), .ZN(p8_mult_21_n352) );
  INV_X1 p8_mult_21_U699 ( .A(p8_mult_21_n167), .ZN(p8_mult_21_n168) );
  INV_X1 p8_mult_21_U708 ( .A(p8_mult_21_n790), .ZN(p8_mult_21_n686) );
  INV_X1 p8_mult_21_U709 ( .A(p8_mult_21_n792), .ZN(p8_mult_21_n685) );
  INV_X1 p8_mult_21_U630 ( .A(p8_mult_21_n788), .ZN(p8_mult_21_n338) );
  INV_X1 p8_mult_21_U656 ( .A(p8_mult_21_n805), .ZN(p8_mult_21_n804) );
  NAND2_X1 p8_mult_21_U695 ( .A1(p8_mult_21_n756), .A2(p8_mult_21_n821), .ZN(
        p8_mult_21_n758) );
  NAND2_X1 p8_mult_21_U702 ( .A1(p8_mult_21_n773), .A2(p8_mult_21_n822), .ZN(
        p8_mult_21_n775) );
  NAND2_X1 p8_mult_21_U710 ( .A1(p8_mult_21_n790), .A2(p8_mult_21_n823), .ZN(
        p8_mult_21_n792) );
  NAND2_X1 p8_mult_21_U723 ( .A1(p8_mult_21_n706), .A2(p8_mult_21_n837), .ZN(
        p8_mult_21_n705) );
  OAI22_X1 p8_mult_21_U493 ( .A1(p8_mult_21_n697), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n698), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n412) );
  NOR2_X1 p8_mult_21_U608 ( .A1(p8_mult_21_n721), .A2(p8_mult_21_n773), .ZN(
        p8_mult_21_n351) );
  OAI22_X1 p8_mult_21_U561 ( .A1(p8_mult_21_n744), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n745), .ZN(p8_mult_21_n375) );
  OAI22_X1 p8_mult_21_U518 ( .A1(p8_mult_21_n713), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n714), .ZN(p8_mult_21_n399) );
  OAI22_X1 p8_mult_21_U584 ( .A1(p8_mult_21_n759), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n760), .ZN(p8_mult_21_n363) );
  OAI22_X1 p8_mult_21_U491 ( .A1(p8_mult_21_n696), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n697), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n413) );
  XNOR2_X1 p8_mult_21_U494 ( .A(B2[9]), .B(reg3_reg[1]), .ZN(p8_mult_21_n697)
         );
  XNOR2_X1 p8_mult_21_U585 ( .A(B2[1]), .B(reg3_reg[9]), .ZN(p8_mult_21_n759)
         );
  OAI22_X1 p8_mult_21_U516 ( .A1(p8_mult_21_n712), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n713), .ZN(p8_mult_21_n400) );
  XNOR2_X1 p8_mult_21_U542 ( .A(B2[5]), .B(reg3_reg[5]), .ZN(p8_mult_21_n729)
         );
  OAI22_X1 p8_mult_21_U559 ( .A1(p8_mult_21_n743), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n744), .ZN(p8_mult_21_n376) );
  XNOR2_X1 p8_mult_21_U562 ( .A(B2[3]), .B(reg3_reg[7]), .ZN(p8_mult_21_n744)
         );
  OAI22_X1 p8_mult_21_U514 ( .A1(p8_mult_21_n711), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n712), .ZN(p8_mult_21_n401) );
  OAI22_X1 p8_mult_21_U557 ( .A1(p8_mult_21_n742), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n743), .ZN(p8_mult_21_n377) );
  XNOR2_X1 p8_mult_21_U560 ( .A(B2[2]), .B(reg3_reg[7]), .ZN(p8_mult_21_n743)
         );
  OAI22_X1 p8_mult_21_U489 ( .A1(p8_mult_21_n695), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n696), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n414) );
  XNOR2_X1 p8_mult_21_U492 ( .A(B2[8]), .B(reg3_reg[1]), .ZN(p8_mult_21_n696)
         );
  NOR2_X1 p8_mult_21_U581 ( .A1(p8_mult_21_n721), .A2(p8_mult_21_n756), .ZN(
        p8_mult_21_n365) );
  XNOR2_X1 p8_mult_21_U540 ( .A(B2[4]), .B(reg3_reg[5]), .ZN(p8_mult_21_n728)
         );
  OAI22_X1 p8_mult_21_U512 ( .A1(p8_mult_21_n710), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n711), .ZN(p8_mult_21_n402) );
  OAI22_X1 p8_mult_21_U487 ( .A1(p8_mult_21_n694), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n695), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n415) );
  XNOR2_X1 p8_mult_21_U490 ( .A(B2[7]), .B(reg3_reg[1]), .ZN(p8_mult_21_n695)
         );
  XNOR2_X1 p8_mult_21_U538 ( .A(B2[3]), .B(reg3_reg[5]), .ZN(p8_mult_21_n727)
         );
  XNOR2_X1 p8_mult_21_U558 ( .A(B2[1]), .B(reg3_reg[7]), .ZN(p8_mult_21_n742)
         );
  OAI22_X1 p8_mult_21_U510 ( .A1(p8_mult_21_n709), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n710), .ZN(p8_mult_21_n403) );
  NOR2_X1 p8_mult_21_U554 ( .A1(p8_mult_21_n721), .A2(p8_mult_21_n739), .ZN(
        p8_mult_21_n379) );
  OAI22_X1 p8_mult_21_U485 ( .A1(p8_mult_21_n693), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n694), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n416) );
  XNOR2_X1 p8_mult_21_U488 ( .A(B2[6]), .B(reg3_reg[1]), .ZN(p8_mult_21_n694)
         );
  XNOR2_X1 p8_mult_21_U536 ( .A(B2[2]), .B(reg3_reg[5]), .ZN(p8_mult_21_n726)
         );
  XNOR2_X1 p8_mult_21_U534 ( .A(B2[1]), .B(reg3_reg[5]), .ZN(p8_mult_21_n725)
         );
  OAI22_X1 p8_mult_21_U483 ( .A1(p8_mult_21_n692), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n693), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n417) );
  XNOR2_X1 p8_mult_21_U486 ( .A(B2[5]), .B(reg3_reg[1]), .ZN(p8_mult_21_n693)
         );
  OAI22_X1 p8_mult_21_U508 ( .A1(p8_mult_21_n708), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n709), .ZN(p8_mult_21_n404) );
  NOR2_X1 p8_mult_21_U422 ( .A1(p8_mult_21_n681), .A2(p8_mult_21_n682), .ZN(
        p8_mult_21_n645) );
  NOR2_X1 p8_mult_21_U420 ( .A1(p8_mult_21_n832), .A2(p8_mult_21_n682), .ZN(
        p8_mult_21_n643) );
  OAI22_X1 p8_mult_21_U506 ( .A1(p8_mult_21_n707), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n708), .ZN(p8_mult_21_n405) );
  OAI22_X1 p8_mult_21_U481 ( .A1(p8_mult_21_n690), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n692), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n418) );
  XNOR2_X1 p8_mult_21_U484 ( .A(B2[4]), .B(reg3_reg[1]), .ZN(p8_mult_21_n692)
         );
  OAI22_X1 p8_mult_21_U480 ( .A1(p8_mult_21_n688), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n690), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n419) );
  XNOR2_X1 p8_mult_21_U482 ( .A(B2[3]), .B(reg3_reg[1]), .ZN(p8_mult_21_n690)
         );
  XNOR2_X1 p8_mult_21_U732 ( .A(B2[2]), .B(reg3_reg[1]), .ZN(p8_mult_21_n688)
         );
  OAI22_X1 p8_mult_21_U520 ( .A1(p8_mult_21_n714), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n715), .ZN(p8_mult_21_n398) );
  OAI22_X1 p8_mult_21_U563 ( .A1(p8_mult_21_n745), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n746), .ZN(p8_mult_21_n374) );
  XNOR2_X1 p8_mult_21_U564 ( .A(B2[4]), .B(reg3_reg[7]), .ZN(p8_mult_21_n745)
         );
  OAI22_X1 p8_mult_21_U495 ( .A1(p8_mult_21_n698), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n699), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n411) );
  XNOR2_X1 p8_mult_21_U496 ( .A(B2[10]), .B(reg3_reg[1]), .ZN(p8_mult_21_n698)
         );
  XNOR2_X1 p8_mult_21_U544 ( .A(B2[6]), .B(reg3_reg[5]), .ZN(p8_mult_21_n730)
         );
  OAI22_X1 p8_mult_21_U586 ( .A1(p8_mult_21_n760), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n761), .ZN(p8_mult_21_n362) );
  XNOR2_X1 p8_mult_21_U587 ( .A(B2[2]), .B(reg3_reg[9]), .ZN(p8_mult_21_n760)
         );
  XNOR2_X1 p8_mult_21_U546 ( .A(B2[7]), .B(reg3_reg[5]), .ZN(p8_mult_21_n731)
         );
  OAI22_X1 p8_mult_21_U565 ( .A1(p8_mult_21_n746), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n747), .ZN(p8_mult_21_n373) );
  XNOR2_X1 p8_mult_21_U566 ( .A(B2[5]), .B(reg3_reg[7]), .ZN(p8_mult_21_n746)
         );
  OAI22_X1 p8_mult_21_U522 ( .A1(p8_mult_21_n715), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n716), .ZN(p8_mult_21_n397) );
  OAI22_X1 p8_mult_21_U611 ( .A1(p8_mult_21_n776), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n777), .ZN(p8_mult_21_n349) );
  XNOR2_X1 p8_mult_21_U612 ( .A(B2[1]), .B(reg3_reg[11]), .ZN(p8_mult_21_n776)
         );
  OAI22_X1 p8_mult_21_U497 ( .A1(p8_mult_21_n699), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n700), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n410) );
  XNOR2_X1 p8_mult_21_U498 ( .A(B2[11]), .B(reg3_reg[1]), .ZN(p8_mult_21_n699)
         );
  NOR2_X1 p8_mult_21_U632 ( .A1(p8_mult_21_n721), .A2(p8_mult_21_n790), .ZN(
        p8_mult_21_n337) );
  OAI22_X1 p8_mult_21_U588 ( .A1(p8_mult_21_n761), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n762), .ZN(p8_mult_21_n361) );
  XNOR2_X1 p8_mult_21_U589 ( .A(B2[3]), .B(reg3_reg[9]), .ZN(p8_mult_21_n761)
         );
  OAI22_X1 p8_mult_21_U590 ( .A1(p8_mult_21_n762), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n763), .ZN(p8_mult_21_n360) );
  XNOR2_X1 p8_mult_21_U591 ( .A(B2[4]), .B(reg3_reg[9]), .ZN(p8_mult_21_n762)
         );
  XNOR2_X1 p8_mult_21_U548 ( .A(B2[8]), .B(reg3_reg[5]), .ZN(p8_mult_21_n732)
         );
  OAI22_X1 p8_mult_21_U613 ( .A1(p8_mult_21_n777), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n778), .ZN(p8_mult_21_n348) );
  XNOR2_X1 p8_mult_21_U614 ( .A(B2[2]), .B(reg3_reg[11]), .ZN(p8_mult_21_n777)
         );
  XNOR2_X1 p8_mult_21_U668 ( .A(p8_mult_21_n816), .B(p8_mult_21_n817), .ZN(
        p8_mult_21_n244) );
  OAI22_X1 p8_mult_21_U524 ( .A1(p8_mult_21_n716), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n717), .ZN(p8_mult_21_n396) );
  OAI22_X1 p8_mult_21_U567 ( .A1(p8_mult_21_n747), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n748), .ZN(p8_mult_21_n372) );
  XNOR2_X1 p8_mult_21_U568 ( .A(B2[6]), .B(reg3_reg[7]), .ZN(p8_mult_21_n747)
         );
  OAI22_X1 p8_mult_21_U499 ( .A1(p8_mult_21_n700), .A2(p8_mult_21_n689), .B1(
        p8_mult_21_n701), .B2(p8_mult_21_n691), .ZN(p8_mult_21_n409) );
  XNOR2_X1 p8_mult_21_U500 ( .A(B2[12]), .B(reg3_reg[1]), .ZN(p8_mult_21_n700)
         );
  OAI22_X1 p8_mult_21_U633 ( .A1(p8_mult_21_n791), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n793), .ZN(p8_mult_21_n336) );
  XNOR2_X1 p8_mult_21_U634 ( .A(reg3_reg[13]), .B(B2[0]), .ZN(p8_mult_21_n791)
         );
  OAI21_X1 p8_mult_21_U666 ( .B1(p8_mult_21_n814), .B2(p8_mult_21_n792), .A(
        p8_mult_21_n815), .ZN(p8_mult_21_n317) );
  OAI22_X1 p8_mult_21_U569 ( .A1(p8_mult_21_n748), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n749), .ZN(p8_mult_21_n371) );
  XNOR2_X1 p8_mult_21_U570 ( .A(B2[7]), .B(reg3_reg[7]), .ZN(p8_mult_21_n748)
         );
  OAI22_X1 p8_mult_21_U635 ( .A1(p8_mult_21_n793), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n794), .ZN(p8_mult_21_n335) );
  XNOR2_X1 p8_mult_21_U636 ( .A(B2[1]), .B(reg3_reg[13]), .ZN(p8_mult_21_n793)
         );
  XNOR2_X1 p8_mult_21_U672 ( .A(B2[9]), .B(reg3_reg[5]), .ZN(p8_mult_21_n733)
         );
  OAI22_X1 p8_mult_21_U673 ( .A1(p8_mult_21_n778), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n779), .ZN(p8_mult_21_n816) );
  XNOR2_X1 p8_mult_21_U675 ( .A(B2[3]), .B(reg3_reg[11]), .ZN(p8_mult_21_n778)
         );
  AOI21_X1 p8_mult_21_U502 ( .B1(p8_mult_21_n689), .B2(p8_mult_21_n691), .A(
        p8_mult_21_n701), .ZN(p8_mult_21_n702) );
  NAND2_X1 p8_mult_21_U733 ( .A1(reg3_reg[1]), .A2(p8_mult_21_n691), .ZN(
        p8_mult_21_n689) );
  OAI22_X1 p8_mult_21_U592 ( .A1(p8_mult_21_n763), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n764), .ZN(p8_mult_21_n359) );
  XNOR2_X1 p8_mult_21_U593 ( .A(B2[5]), .B(reg3_reg[9]), .ZN(p8_mult_21_n763)
         );
  OAI22_X1 p8_mult_21_U526 ( .A1(p8_mult_21_n717), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n718), .ZN(p8_mult_21_n395) );
  AOI21_X1 p8_mult_21_U529 ( .B1(p8_mult_21_n705), .B2(p8_mult_21_n706), .A(
        p8_mult_21_n720), .ZN(p8_mult_21_n719) );
  OAI22_X1 p8_mult_21_U639 ( .A1(p8_mult_21_n795), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n796), .ZN(p8_mult_21_n333) );
  OAI22_X1 p8_mult_21_U598 ( .A1(p8_mult_21_n766), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n767), .ZN(p8_mult_21_n356) );
  OAI22_X1 p8_mult_21_U641 ( .A1(p8_mult_21_n796), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n797), .ZN(p8_mult_21_n332) );
  XNOR2_X1 p8_mult_21_U642 ( .A(B2[4]), .B(reg3_reg[13]), .ZN(p8_mult_21_n796)
         );
  OAI22_X1 p8_mult_21_U594 ( .A1(p8_mult_21_n764), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n765), .ZN(p8_mult_21_n358) );
  XNOR2_X1 p8_mult_21_U595 ( .A(B2[6]), .B(reg3_reg[9]), .ZN(p8_mult_21_n764)
         );
  OAI22_X1 p8_mult_21_U571 ( .A1(p8_mult_21_n749), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n750), .ZN(p8_mult_21_n370) );
  XNOR2_X1 p8_mult_21_U572 ( .A(B2[8]), .B(reg3_reg[7]), .ZN(p8_mult_21_n749)
         );
  OAI22_X1 p8_mult_21_U637 ( .A1(p8_mult_21_n794), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n795), .ZN(p8_mult_21_n334) );
  XNOR2_X1 p8_mult_21_U640 ( .A(B2[3]), .B(reg3_reg[13]), .ZN(p8_mult_21_n795)
         );
  XNOR2_X1 p8_mult_21_U638 ( .A(B2[2]), .B(reg3_reg[13]), .ZN(p8_mult_21_n794)
         );
  OAI22_X1 p8_mult_21_U573 ( .A1(p8_mult_21_n750), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n751), .ZN(p8_mult_21_n369) );
  XNOR2_X1 p8_mult_21_U574 ( .A(B2[9]), .B(reg3_reg[7]), .ZN(p8_mult_21_n750)
         );
  OAI22_X1 p8_mult_21_U677 ( .A1(p8_mult_21_n718), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n720), .ZN(p8_mult_21_n231) );
  XNOR2_X1 p8_mult_21_U724 ( .A(p8_mult_21_n819), .B(reg3_reg[2]), .ZN(
        p8_mult_21_n837) );
  OAI22_X1 p8_mult_21_U615 ( .A1(p8_mult_21_n779), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n780), .ZN(p8_mult_21_n346) );
  XNOR2_X1 p8_mult_21_U674 ( .A(B2[4]), .B(reg3_reg[11]), .ZN(p8_mult_21_n779)
         );
  XNOR2_X1 p8_mult_21_U671 ( .A(B2[10]), .B(reg3_reg[5]), .ZN(p8_mult_21_n734)
         );
  OAI22_X1 p8_mult_21_U596 ( .A1(p8_mult_21_n765), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n766), .ZN(p8_mult_21_n357) );
  XNOR2_X1 p8_mult_21_U599 ( .A(B2[8]), .B(reg3_reg[9]), .ZN(p8_mult_21_n766)
         );
  XNOR2_X1 p8_mult_21_U597 ( .A(B2[7]), .B(reg3_reg[9]), .ZN(p8_mult_21_n765)
         );
  XNOR2_X1 p8_mult_21_U551 ( .A(B2[11]), .B(reg3_reg[5]), .ZN(p8_mult_21_n735)
         );
  OAI22_X1 p8_mult_21_U616 ( .A1(p8_mult_21_n780), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n781), .ZN(p8_mult_21_n345) );
  XNOR2_X1 p8_mult_21_U617 ( .A(B2[5]), .B(reg3_reg[11]), .ZN(p8_mult_21_n780)
         );
  OAI22_X1 p8_mult_21_U618 ( .A1(p8_mult_21_n781), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n782), .ZN(p8_mult_21_n344) );
  XNOR2_X1 p8_mult_21_U619 ( .A(B2[6]), .B(reg3_reg[11]), .ZN(p8_mult_21_n781)
         );
  OAI22_X1 p8_mult_21_U575 ( .A1(p8_mult_21_n751), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n752), .ZN(p8_mult_21_n368) );
  XNOR2_X1 p8_mult_21_U576 ( .A(B2[10]), .B(reg3_reg[7]), .ZN(p8_mult_21_n751)
         );
  OAI22_X1 p8_mult_21_U577 ( .A1(p8_mult_21_n752), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n753), .ZN(p8_mult_21_n367) );
  XNOR2_X1 p8_mult_21_U578 ( .A(B2[11]), .B(reg3_reg[7]), .ZN(p8_mult_21_n752)
         );
  OAI22_X1 p8_mult_21_U620 ( .A1(p8_mult_21_n782), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n783), .ZN(p8_mult_21_n343) );
  XNOR2_X1 p8_mult_21_U621 ( .A(B2[7]), .B(reg3_reg[11]), .ZN(p8_mult_21_n782)
         );
  OAI22_X1 p8_mult_21_U600 ( .A1(p8_mult_21_n767), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n768), .ZN(p8_mult_21_n355) );
  XNOR2_X1 p8_mult_21_U601 ( .A(B2[9]), .B(reg3_reg[9]), .ZN(p8_mult_21_n767)
         );
  OAI22_X1 p8_mult_21_U602 ( .A1(p8_mult_21_n768), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n769), .ZN(p8_mult_21_n354) );
  XNOR2_X1 p8_mult_21_U603 ( .A(B2[10]), .B(reg3_reg[9]), .ZN(p8_mult_21_n768)
         );
  OAI22_X1 p8_mult_21_U643 ( .A1(p8_mult_21_n797), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n798), .ZN(p8_mult_21_n331) );
  XNOR2_X1 p8_mult_21_U644 ( .A(B2[5]), .B(reg3_reg[13]), .ZN(p8_mult_21_n797)
         );
  XNOR2_X1 p8_mult_21_U682 ( .A(B2[13]), .B(reg3_reg[5]), .ZN(p8_mult_21_n738)
         );
  XNOR2_X1 p8_mult_21_U683 ( .A(p8_mult_21_n806), .B(reg3_reg[4]), .ZN(
        p8_mult_21_n818) );
  XNOR2_X1 p8_mult_21_U684 ( .A(B2[12]), .B(reg3_reg[5]), .ZN(p8_mult_21_n736)
         );
  OAI22_X1 p8_mult_21_U622 ( .A1(p8_mult_21_n783), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n784), .ZN(p8_mult_21_n342) );
  XNOR2_X1 p8_mult_21_U623 ( .A(B2[8]), .B(reg3_reg[11]), .ZN(p8_mult_21_n783)
         );
  OAI22_X1 p8_mult_21_U645 ( .A1(p8_mult_21_n798), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n799), .ZN(p8_mult_21_n330) );
  XNOR2_X1 p8_mult_21_U646 ( .A(B2[6]), .B(reg3_reg[13]), .ZN(p8_mult_21_n798)
         );
  OAI22_X1 p8_mult_21_U604 ( .A1(p8_mult_21_n769), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n770), .ZN(p8_mult_21_n353) );
  XNOR2_X1 p8_mult_21_U605 ( .A(B2[11]), .B(reg3_reg[9]), .ZN(p8_mult_21_n769)
         );
  OAI22_X1 p8_mult_21_U624 ( .A1(p8_mult_21_n784), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n785), .ZN(p8_mult_21_n341) );
  XNOR2_X1 p8_mult_21_U625 ( .A(B2[9]), .B(reg3_reg[11]), .ZN(p8_mult_21_n784)
         );
  AOI21_X1 p8_mult_21_U580 ( .B1(p8_mult_21_n741), .B2(p8_mult_21_n739), .A(
        p8_mult_21_n755), .ZN(p8_mult_21_n754) );
  OAI22_X1 p8_mult_21_U647 ( .A1(p8_mult_21_n799), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n800), .ZN(p8_mult_21_n329) );
  XNOR2_X1 p8_mult_21_U648 ( .A(B2[7]), .B(reg3_reg[13]), .ZN(p8_mult_21_n799)
         );
  OAI22_X1 p8_mult_21_U686 ( .A1(p8_mult_21_n753), .A2(p8_mult_21_n741), .B1(
        p8_mult_21_n739), .B2(p8_mult_21_n755), .ZN(p8_mult_21_n191) );
  XNOR2_X1 p8_mult_21_U687 ( .A(B2[13]), .B(reg3_reg[7]), .ZN(p8_mult_21_n755)
         );
  XNOR2_X1 p8_mult_21_U689 ( .A(p8_mult_21_n808), .B(reg3_reg[6]), .ZN(
        p8_mult_21_n820) );
  XNOR2_X1 p8_mult_21_U691 ( .A(B2[12]), .B(reg3_reg[7]), .ZN(p8_mult_21_n753)
         );
  OAI22_X1 p8_mult_21_U628 ( .A1(p8_mult_21_n786), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n787), .ZN(p8_mult_21_n339) );
  OAI22_X1 p8_mult_21_U626 ( .A1(p8_mult_21_n785), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n786), .ZN(p8_mult_21_n340) );
  XNOR2_X1 p8_mult_21_U629 ( .A(B2[11]), .B(reg3_reg[11]), .ZN(p8_mult_21_n786) );
  XNOR2_X1 p8_mult_21_U627 ( .A(B2[10]), .B(reg3_reg[11]), .ZN(p8_mult_21_n785) );
  OAI22_X1 p8_mult_21_U649 ( .A1(p8_mult_21_n800), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n801), .ZN(p8_mult_21_n328) );
  XNOR2_X1 p8_mult_21_U650 ( .A(B2[8]), .B(reg3_reg[13]), .ZN(p8_mult_21_n800)
         );
  AOI21_X1 p8_mult_21_U607 ( .B1(p8_mult_21_n758), .B2(p8_mult_21_n756), .A(
        p8_mult_21_n772), .ZN(p8_mult_21_n771) );
  OAI22_X1 p8_mult_21_U693 ( .A1(p8_mult_21_n770), .A2(p8_mult_21_n758), .B1(
        p8_mult_21_n756), .B2(p8_mult_21_n772), .ZN(p8_mult_21_n177) );
  XNOR2_X1 p8_mult_21_U694 ( .A(B2[13]), .B(reg3_reg[9]), .ZN(p8_mult_21_n772)
         );
  XNOR2_X1 p8_mult_21_U696 ( .A(p8_mult_21_n810), .B(reg3_reg[8]), .ZN(
        p8_mult_21_n821) );
  XNOR2_X1 p8_mult_21_U698 ( .A(B2[12]), .B(reg3_reg[9]), .ZN(p8_mult_21_n770)
         );
  OAI22_X1 p8_mult_21_U651 ( .A1(p8_mult_21_n801), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n802), .ZN(p8_mult_21_n327) );
  XNOR2_X1 p8_mult_21_U652 ( .A(B2[9]), .B(reg3_reg[13]), .ZN(p8_mult_21_n801)
         );
  OAI22_X1 p8_mult_21_U653 ( .A1(p8_mult_21_n802), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n803), .ZN(p8_mult_21_n326) );
  XNOR2_X1 p8_mult_21_U654 ( .A(B2[10]), .B(reg3_reg[13]), .ZN(p8_mult_21_n802) );
  AOI22_X1 p8_mult_21_U706 ( .A1(p8_mult_21_n805), .A2(p8_mult_21_n685), .B1(
        p8_mult_21_n686), .B2(p8_mult_21_n687), .ZN(p8_mult_21_n162) );
  XNOR2_X1 p8_mult_21_U707 ( .A(B2[13]), .B(p8_mult_21_n814), .ZN(
        p8_mult_21_n687) );
  AOI21_X1 p8_mult_21_U631 ( .B1(p8_mult_21_n775), .B2(p8_mult_21_n773), .A(
        p8_mult_21_n789), .ZN(p8_mult_21_n788) );
  OAI22_X1 p8_mult_21_U700 ( .A1(p8_mult_21_n787), .A2(p8_mult_21_n775), .B1(
        p8_mult_21_n773), .B2(p8_mult_21_n789), .ZN(p8_mult_21_n167) );
  XNOR2_X1 p8_mult_21_U701 ( .A(B2[13]), .B(reg3_reg[11]), .ZN(p8_mult_21_n789) );
  XNOR2_X1 p8_mult_21_U703 ( .A(p8_mult_21_n812), .B(reg3_reg[10]), .ZN(
        p8_mult_21_n822) );
  XNOR2_X1 p8_mult_21_U705 ( .A(B2[12]), .B(reg3_reg[11]), .ZN(p8_mult_21_n787) );
  OAI22_X1 p8_mult_21_U655 ( .A1(p8_mult_21_n803), .A2(p8_mult_21_n792), .B1(
        p8_mult_21_n790), .B2(p8_mult_21_n804), .ZN(p8_mult_21_n325) );
  XNOR2_X1 p8_mult_21_U711 ( .A(p8_mult_21_n814), .B(reg3_reg[12]), .ZN(
        p8_mult_21_n823) );
  XNOR2_X1 p8_mult_21_U657 ( .A(B2[11]), .B(reg3_reg[13]), .ZN(p8_mult_21_n803) );
  XOR2_X1 p8_mult_21_U737 ( .A(reg3_reg[2]), .B(reg3_reg[1]), .Z(
        p8_mult_21_n836) );
  XOR2_X1 p8_mult_21_U714 ( .A(B2[12]), .B(reg3_reg[13]), .Z(p8_mult_21_n805)
         );
  NAND3_X1 p8_mult_21_U667 ( .A1(p8_mult_21_n686), .A2(p8_mult_21_n721), .A3(
        reg3_reg[13]), .ZN(p8_mult_21_n815) );
  XOR2_X1 p8_mult_21_U503 ( .A(B2[13]), .B(p8_mult_21_n703), .Z(
        p8_mult_21_n701) );
  XOR2_X1 p8_mult_21_U460 ( .A(p8_mult_21_n657), .B(p8_mult_21_n670), .Z(
        temp3[0]) );
  XOR2_X1 p8_mult_21_U459 ( .A(p8_mult_21_n246), .B(p8_mult_21_n257), .Z(
        p8_mult_21_n670) );
  XOR2_X1 p8_mult_21_U454 ( .A(p8_mult_21_n148), .B(p8_mult_21_n666), .Z(
        temp3[1]) );
  XOR2_X1 p8_mult_21_U453 ( .A(p8_mult_21_n234), .B(p8_mult_21_n245), .Z(
        p8_mult_21_n666) );
  XOR2_X1 p8_mult_21_U434 ( .A(p8_mult_21_n147), .B(p8_mult_21_n650), .Z(
        temp3[2]) );
  XOR2_X1 p8_mult_21_U433 ( .A(p8_mult_21_n222), .B(p8_mult_21_n233), .Z(
        p8_mult_21_n650) );
  XOR2_X1 p8_mult_21_U428 ( .A(p8_mult_21_n143), .B(p8_mult_21_n646), .Z(
        temp3[6]) );
  XOR2_X1 p8_mult_21_U427 ( .A(p8_mult_21_n193), .B(p8_mult_21_n186), .Z(
        p8_mult_21_n646) );
  HA_X1 p8_mult_21_U145 ( .A(p8_mult_21_n406), .B(p8_mult_21_n419), .CO(
        p8_mult_21_n315), .S(p8_mult_21_n316) );
  FA_X1 p8_mult_21_U144 ( .A(p8_mult_21_n418), .B(p8_mult_21_n393), .CI(
        p8_mult_21_n405), .CO(p8_mult_21_n313), .S(p8_mult_21_n314) );
  FA_X1 p8_mult_21_U141 ( .A(p8_mult_21_n416), .B(p8_mult_21_n379), .CI(
        p8_mult_21_n403), .CO(p8_mult_21_n307), .S(p8_mult_21_n308) );
  FA_X1 p8_mult_21_U138 ( .A(p8_mult_21_n390), .B(p8_mult_21_n415), .CI(
        p8_mult_21_n402), .CO(p8_mult_21_n301), .S(p8_mult_21_n302) );
  FA_X1 p8_mult_21_U137 ( .A(p8_mult_21_n307), .B(p8_mult_21_n304), .CI(
        p8_mult_21_n302), .CO(p8_mult_21_n299), .S(p8_mult_21_n300) );
  FA_X1 p8_mult_21_U136 ( .A(p8_mult_21_n389), .B(p8_mult_21_n365), .CI(
        p8_mult_21_n414), .CO(p8_mult_21_n297), .S(p8_mult_21_n298) );
  FA_X1 p8_mult_21_U135 ( .A(p8_mult_21_n377), .B(p8_mult_21_n401), .CI(
        p8_mult_21_n303), .CO(p8_mult_21_n295), .S(p8_mult_21_n296) );
  FA_X1 p8_mult_21_U134 ( .A(p8_mult_21_n298), .B(p8_mult_21_n301), .CI(
        p8_mult_21_n296), .CO(p8_mult_21_n293), .S(p8_mult_21_n294) );
  FA_X1 p8_mult_21_U132 ( .A(p8_mult_21_n376), .B(p8_mult_21_n388), .CI(
        p8_mult_21_n400), .CO(p8_mult_21_n289), .S(p8_mult_21_n290) );
  FA_X1 p8_mult_21_U129 ( .A(p8_mult_21_n375), .B(p8_mult_21_n351), .CI(
        p8_mult_21_n412), .CO(p8_mult_21_n283), .S(p8_mult_21_n284) );
  FA_X1 p8_mult_21_U128 ( .A(p8_mult_21_n363), .B(p8_mult_21_n399), .CI(
        p8_mult_21_n387), .CO(p8_mult_21_n281), .S(p8_mult_21_n282) );
  FA_X1 p8_mult_21_U127 ( .A(p8_mult_21_n289), .B(p8_mult_21_n291), .CI(
        p8_mult_21_n284), .CO(p8_mult_21_n279), .S(p8_mult_21_n280) );
  FA_X1 p8_mult_21_U124 ( .A(p8_mult_21_n362), .B(p8_mult_21_n386), .CI(
        p8_mult_21_n411), .CO(p8_mult_21_n273), .S(p8_mult_21_n274) );
  FA_X1 p8_mult_21_U123 ( .A(p8_mult_21_n374), .B(p8_mult_21_n398), .CI(
        p8_mult_21_n276), .CO(p8_mult_21_n271), .S(p8_mult_21_n272) );
  FA_X1 p8_mult_21_U122 ( .A(p8_mult_21_n281), .B(p8_mult_21_n283), .CI(
        p8_mult_21_n274), .CO(p8_mult_21_n269), .S(p8_mult_21_n270) );
  FA_X1 p8_mult_21_U121 ( .A(p8_mult_21_n279), .B(p8_mult_21_n272), .CI(
        p8_mult_21_n270), .CO(p8_mult_21_n267), .S(p8_mult_21_n268) );
  FA_X1 p8_mult_21_U120 ( .A(p8_mult_21_n361), .B(p8_mult_21_n337), .CI(
        p8_mult_21_n410), .CO(p8_mult_21_n265), .S(p8_mult_21_n266) );
  FA_X1 p8_mult_21_U109 ( .A(p8_mult_21_n349), .B(p8_mult_21_n397), .CI(
        p8_mult_21_n373), .CO(p8_mult_21_n263), .S(p8_mult_21_n264) );
  FA_X1 p8_mult_21_U108 ( .A(p8_mult_21_n275), .B(p8_mult_21_n385), .CI(
        p8_mult_21_n273), .CO(p8_mult_21_n261), .S(p8_mult_21_n262) );
  FA_X1 p8_mult_21_U107 ( .A(p8_mult_21_n264), .B(p8_mult_21_n266), .CI(
        p8_mult_21_n271), .CO(p8_mult_21_n259), .S(p8_mult_21_n260) );
  FA_X1 p8_mult_21_U106 ( .A(p8_mult_21_n262), .B(p8_mult_21_n269), .CI(
        p8_mult_21_n260), .CO(p8_mult_21_n257), .S(p8_mult_21_n258) );
  HA_X1 p8_mult_21_U105 ( .A(p8_mult_21_n317), .B(p8_mult_21_n336), .CO(
        p8_mult_21_n255), .S(p8_mult_21_n256) );
  FA_X1 p8_mult_21_U104 ( .A(p8_mult_21_n409), .B(p8_mult_21_n372), .CI(
        p8_mult_21_n396), .CO(p8_mult_21_n253), .S(p8_mult_21_n254) );
  FA_X1 p8_mult_21_U103 ( .A(p8_mult_21_n348), .B(p8_mult_21_n384), .CI(
        p8_mult_21_n360), .CO(p8_mult_21_n251), .S(p8_mult_21_n252) );
  FA_X1 p8_mult_21_U102 ( .A(p8_mult_21_n265), .B(p8_mult_21_n256), .CI(
        p8_mult_21_n263), .CO(p8_mult_21_n249), .S(p8_mult_21_n250) );
  FA_X1 p8_mult_21_U101 ( .A(p8_mult_21_n254), .B(p8_mult_21_n252), .CI(
        p8_mult_21_n261), .CO(p8_mult_21_n247), .S(p8_mult_21_n248) );
  FA_X1 p8_mult_21_U100 ( .A(p8_mult_21_n259), .B(p8_mult_21_n250), .CI(
        p8_mult_21_n248), .CO(p8_mult_21_n245), .S(p8_mult_21_n246) );
  FA_X1 p8_mult_21_U97 ( .A(p8_mult_21_n395), .B(p8_mult_21_n359), .CI(
        p8_mult_21_n408), .CO(p8_mult_21_n241), .S(p8_mult_21_n242) );
  FA_X1 p8_mult_21_U96 ( .A(p8_mult_21_n335), .B(p8_mult_21_n371), .CI(
        p8_mult_21_n255), .CO(p8_mult_21_n239), .S(p8_mult_21_n240) );
  FA_X1 p8_mult_21_U95 ( .A(p8_mult_21_n253), .B(p8_mult_21_n244), .CI(
        p8_mult_21_n251), .CO(p8_mult_21_n237), .S(p8_mult_21_n238) );
  FA_X1 p8_mult_21_U94 ( .A(p8_mult_21_n240), .B(p8_mult_21_n242), .CI(
        p8_mult_21_n249), .CO(p8_mult_21_n235), .S(p8_mult_21_n236) );
  FA_X1 p8_mult_21_U93 ( .A(p8_mult_21_n247), .B(p8_mult_21_n238), .CI(
        p8_mult_21_n236), .CO(p8_mult_21_n233), .S(p8_mult_21_n234) );
  FA_X1 p8_mult_21_U91 ( .A(p8_mult_21_n382), .B(p8_mult_21_n346), .CI(
        p8_mult_21_n232), .CO(p8_mult_21_n229), .S(p8_mult_21_n230) );
  FA_X1 p8_mult_21_U90 ( .A(p8_mult_21_n334), .B(p8_mult_21_n370), .CI(
        p8_mult_21_n358), .CO(p8_mult_21_n227), .S(p8_mult_21_n228) );
  FA_X1 p8_mult_21_U89 ( .A(p8_mult_21_n241), .B(p8_mult_21_n243), .CI(
        p8_mult_21_n239), .CO(p8_mult_21_n225), .S(p8_mult_21_n226) );
  FA_X1 p8_mult_21_U88 ( .A(p8_mult_21_n230), .B(p8_mult_21_n228), .CI(
        p8_mult_21_n237), .CO(p8_mult_21_n223), .S(p8_mult_21_n224) );
  FA_X1 p8_mult_21_U87 ( .A(p8_mult_21_n235), .B(p8_mult_21_n226), .CI(
        p8_mult_21_n224), .CO(p8_mult_21_n221), .S(p8_mult_21_n222) );
  FA_X1 p8_mult_21_U86 ( .A(p8_mult_21_n231), .B(p8_mult_21_n333), .CI(
        p8_mult_21_n394), .CO(p8_mult_21_n219), .S(p8_mult_21_n220) );
  FA_X1 p8_mult_21_U85 ( .A(p8_mult_21_n345), .B(p8_mult_21_n381), .CI(
        p8_mult_21_n357), .CO(p8_mult_21_n217), .S(p8_mult_21_n218) );
  FA_X1 p8_mult_21_U84 ( .A(p8_mult_21_n229), .B(p8_mult_21_n369), .CI(
        p8_mult_21_n227), .CO(p8_mult_21_n215), .S(p8_mult_21_n216) );
  FA_X1 p8_mult_21_U83 ( .A(p8_mult_21_n220), .B(p8_mult_21_n218), .CI(
        p8_mult_21_n225), .CO(p8_mult_21_n213), .S(p8_mult_21_n214) );
  FA_X1 p8_mult_21_U82 ( .A(p8_mult_21_n223), .B(p8_mult_21_n216), .CI(
        p8_mult_21_n214), .CO(p8_mult_21_n211), .S(p8_mult_21_n212) );
  FA_X1 p8_mult_21_U80 ( .A(p8_mult_21_n368), .B(p8_mult_21_n344), .CI(
        p8_mult_21_n210), .CO(p8_mult_21_n207), .S(p8_mult_21_n208) );
  FA_X1 p8_mult_21_U79 ( .A(p8_mult_21_n332), .B(p8_mult_21_n356), .CI(
        p8_mult_21_n219), .CO(p8_mult_21_n205), .S(p8_mult_21_n206) );
  FA_X1 p8_mult_21_U78 ( .A(p8_mult_21_n208), .B(p8_mult_21_n217), .CI(
        p8_mult_21_n215), .CO(p8_mult_21_n203), .S(p8_mult_21_n204) );
  FA_X1 p8_mult_21_U77 ( .A(p8_mult_21_n213), .B(p8_mult_21_n206), .CI(
        p8_mult_21_n204), .CO(p8_mult_21_n201), .S(p8_mult_21_n202) );
  FA_X1 p8_mult_21_U76 ( .A(p8_mult_21_n209), .B(p8_mult_21_n331), .CI(
        p8_mult_21_n380), .CO(p8_mult_21_n199), .S(p8_mult_21_n200) );
  FA_X1 p8_mult_21_U75 ( .A(p8_mult_21_n355), .B(p8_mult_21_n343), .CI(
        p8_mult_21_n367), .CO(p8_mult_21_n197), .S(p8_mult_21_n198) );
  FA_X1 p8_mult_21_U74 ( .A(p8_mult_21_n198), .B(p8_mult_21_n207), .CI(
        p8_mult_21_n200), .CO(p8_mult_21_n195), .S(p8_mult_21_n196) );
  FA_X1 p8_mult_21_U73 ( .A(p8_mult_21_n203), .B(p8_mult_21_n205), .CI(
        p8_mult_21_n196), .CO(p8_mult_21_n193), .S(p8_mult_21_n194) );
  FA_X1 p8_mult_21_U71 ( .A(p8_mult_21_n330), .B(p8_mult_21_n342), .CI(
        p8_mult_21_n192), .CO(p8_mult_21_n189), .S(p8_mult_21_n190) );
  FA_X1 p8_mult_21_U70 ( .A(p8_mult_21_n199), .B(p8_mult_21_n354), .CI(
        p8_mult_21_n197), .CO(p8_mult_21_n187), .S(p8_mult_21_n188) );
  FA_X1 p8_mult_21_U69 ( .A(p8_mult_21_n188), .B(p8_mult_21_n190), .CI(
        p8_mult_21_n195), .CO(p8_mult_21_n185), .S(p8_mult_21_n186) );
  FA_X1 p8_mult_21_U68 ( .A(p8_mult_21_n191), .B(p8_mult_21_n329), .CI(
        p8_mult_21_n366), .CO(p8_mult_21_n183), .S(p8_mult_21_n184) );
  FA_X1 p8_mult_21_U67 ( .A(p8_mult_21_n341), .B(p8_mult_21_n353), .CI(
        p8_mult_21_n189), .CO(p8_mult_21_n181), .S(p8_mult_21_n182) );
  FA_X1 p8_mult_21_U66 ( .A(p8_mult_21_n187), .B(p8_mult_21_n184), .CI(
        p8_mult_21_n182), .CO(p8_mult_21_n179), .S(p8_mult_21_n180) );
  FA_X1 p8_mult_21_U64 ( .A(p8_mult_21_n328), .B(p8_mult_21_n340), .CI(
        p8_mult_21_n178), .CO(p8_mult_21_n175), .S(p8_mult_21_n176) );
  FA_X1 p8_mult_21_U63 ( .A(p8_mult_21_n176), .B(p8_mult_21_n183), .CI(
        p8_mult_21_n181), .CO(p8_mult_21_n173), .S(p8_mult_21_n174) );
  FA_X1 p8_mult_21_U62 ( .A(p8_mult_21_n327), .B(p8_mult_21_n177), .CI(
        p8_mult_21_n352), .CO(p8_mult_21_n171), .S(p8_mult_21_n172) );
  FA_X1 p8_mult_21_U61 ( .A(p8_mult_21_n175), .B(p8_mult_21_n339), .CI(
        p8_mult_21_n172), .CO(p8_mult_21_n169), .S(p8_mult_21_n170) );
  FA_X1 p8_mult_21_U59 ( .A(p8_mult_21_n168), .B(p8_mult_21_n326), .CI(
        p8_mult_21_n171), .CO(p8_mult_21_n165), .S(p8_mult_21_n166) );
  FA_X1 p8_mult_21_U58 ( .A(p8_mult_21_n325), .B(p8_mult_21_n167), .CI(
        p8_mult_21_n338), .CO(p8_mult_21_n163), .S(p8_mult_21_n164) );
  FA_X1 p8_mult_21_U41 ( .A(p8_mult_21_n212), .B(p8_mult_21_n221), .CI(
        p8_mult_21_n146), .CO(p8_mult_21_n145), .S(temp3[3]) );
  FA_X1 p8_mult_21_U40 ( .A(p8_mult_21_n202), .B(p8_mult_21_n211), .CI(
        p8_mult_21_n145), .CO(p8_mult_21_n144), .S(temp3[4]) );
  FA_X1 p8_mult_21_U39 ( .A(p8_mult_21_n194), .B(p8_mult_21_n201), .CI(
        p8_mult_21_n144), .CO(p8_mult_21_n143), .S(temp3[5]) );
  FA_X1 p8_mult_21_U37 ( .A(p8_mult_21_n180), .B(p8_mult_21_n185), .CI(
        p8_mult_21_n142), .CO(p8_mult_21_n141), .S(temp3[7]) );
  FA_X1 p8_mult_21_U30 ( .A(p8_mult_21_n174), .B(p8_mult_21_n179), .CI(
        p8_mult_21_n141), .CO(p8_mult_21_n140), .S(temp3[8]) );
  FA_X1 p8_mult_21_U20 ( .A(p8_mult_21_n170), .B(p8_mult_21_n173), .CI(
        p8_mult_21_n140), .CO(p8_mult_21_n139), .S(temp3[9]) );
  FA_X1 p8_mult_21_U10 ( .A(p8_mult_21_n166), .B(p8_mult_21_n169), .CI(
        p8_mult_21_n139), .CO(p8_mult_21_n138), .S(temp3[10]) );
  FA_X1 p8_mult_21_U9 ( .A(p8_mult_21_n165), .B(p8_mult_21_n164), .CI(
        p8_mult_21_n138), .CO(p8_mult_21_n137), .S(temp3[11]) );
  FA_X1 p8_mult_21_U8 ( .A(p8_mult_21_n163), .B(p8_mult_21_n162), .CI(
        p8_mult_21_n137), .CO(p8_mult_21_n136), .S(temp3[12]) );
  INV_X1 p9_mult_21_U438 ( .A(p9_mult_21_n875), .ZN(p9_mult_21_n873) );
  INV_X1 p9_mult_21_U463 ( .A(p9_mult_21_n915), .ZN(p9_mult_21_n914) );
  INV_X1 p9_mult_21_U484 ( .A(p9_mult_21_n947), .ZN(p9_mult_21_n945) );
  INV_X1 p9_mult_21_U494 ( .A(p9_mult_21_n963), .ZN(p9_mult_21_n962) );
  INV_X1 p9_mult_21_U496 ( .A(p9_mult_21_n966), .ZN(p9_mult_21_n965) );
  INV_X1 p9_mult_21_U837 ( .A(p9_mult_21_n1352), .ZN(p9_mult_21_n1387) );
  INV_X1 p9_mult_21_U652 ( .A(p9_mult_21_n1194), .ZN(p9_mult_21_n1191) );
  INV_X1 p9_mult_21_U750 ( .A(p9_mult_21_n1330), .ZN(p9_mult_21_n1201) );
  INV_X1 p9_mult_21_U661 ( .A(p9_mult_21_n1219), .ZN(p9_mult_21_n1218) );
  INV_X1 p9_mult_21_U709 ( .A(p9_mult_21_n1300), .ZN(p9_mult_21_n1299) );
  INV_X1 p9_mult_21_U418 ( .A(p9_mult_21_n1303), .ZN(p9_mult_21_n845) );
  INV_X1 p9_mult_21_U677 ( .A(p9_mult_21_n1265), .ZN(p9_mult_21_n1262) );
  INV_X1 p9_mult_21_U412 ( .A(p9_mult_21_n1271), .ZN(p9_mult_21_n839) );
  INV_X1 p9_mult_21_U414 ( .A(p9_mult_21_n1286), .ZN(p9_mult_21_n841) );
  INV_X1 p9_mult_21_U763 ( .A(p9_mult_21_n1340), .ZN(p9_mult_21_n1338) );
  INV_X1 p9_mult_21_U726 ( .A(p9_mult_21_n1309), .ZN(p9_mult_21_n1209) );
  INV_X1 p9_mult_21_U745 ( .A(p9_mult_21_n985), .ZN(p9_mult_21_n952) );
  INV_X1 p9_mult_21_U785 ( .A(p9_mult_21_n1362), .ZN(p9_mult_21_n1356) );
  INV_X1 p9_mult_21_U835 ( .A(p9_mult_21_n1386), .ZN(p9_mult_21_n1383) );
  INV_X1 p9_mult_21_U630 ( .A(p9_mult_21_n1158), .ZN(p9_mult_21_n1157) );
  INV_X1 p9_mult_21_U801 ( .A(p9_mult_21_n1360), .ZN(p9_mult_21_n1369) );
  INV_X1 p9_mult_21_U627 ( .A(p9_mult_21_n1151), .ZN(p9_mult_21_n1107) );
  INV_X1 p9_mult_21_U814 ( .A(p9_mult_21_n1167), .ZN(p9_mult_21_n1373) );
  INV_X1 p9_mult_21_U571 ( .A(p9_mult_21_n1070), .ZN(p9_mult_21_n1052) );
  INV_X1 p9_mult_21_U562 ( .A(p9_mult_21_n1059), .ZN(p9_mult_21_n1058) );
  INV_X1 p9_mult_21_U566 ( .A(p9_mult_21_n1061), .ZN(p9_mult_21_n1060) );
  INV_X1 p9_mult_21_U578 ( .A(p9_mult_21_n1084), .ZN(p9_mult_21_n1083) );
  INV_X1 p9_mult_21_U581 ( .A(p9_mult_21_n1086), .ZN(p9_mult_21_n1085) );
  AND2_X1 p9_mult_21_U611 ( .A1(p9_mult_21_n1123), .A2(p9_mult_21_n1124), .ZN(
        p9_mult_21_n1097) );
  INV_X1 p9_mult_21_U869 ( .A(p9_mult_21_n903), .ZN(p9_mult_21_n881) );
  INV_X1 p9_mult_21_U881 ( .A(B3[4]), .ZN(p9_mult_21_n1094) );
  INV_X1 p9_mult_21_U872 ( .A(B3[2]), .ZN(p9_mult_21_n1175) );
  AND2_X1 p9_mult_21_U640 ( .A1(p9_mult_21_n1172), .A2(p9_mult_21_n1173), .ZN(
        p9_mult_21_n1128) );
  INV_X1 p9_mult_21_U519 ( .A(p9_mult_21_n994), .ZN(p9_mult_21_n992) );
  INV_X1 p9_mult_21_U521 ( .A(p9_mult_21_n998), .ZN(p9_mult_21_n995) );
  INV_X1 p9_mult_21_U803 ( .A(p9_mult_21_n1044), .ZN(p9_mult_21_n1022) );
  INV_X1 p9_mult_21_U850 ( .A(B3[5]), .ZN(p9_mult_21_n1062) );
  INV_X1 p9_mult_21_U843 ( .A(B3[8]), .ZN(p9_mult_21_n955) );
  INV_X1 p9_mult_21_U533 ( .A(p9_mult_21_n1016), .ZN(p9_mult_21_n999) );
  INV_X1 p9_mult_21_U535 ( .A(p9_mult_21_n993), .ZN(p9_mult_21_n1019) );
  INV_X1 p9_mult_21_U853 ( .A(B3[6]), .ZN(p9_mult_21_n1025) );
  INV_X1 p9_mult_21_U819 ( .A(B3[7]), .ZN(p9_mult_21_n983) );
  INV_X1 p9_mult_21_U873 ( .A(p9_mult_21_n911), .ZN(p9_mult_21_n880) );
  INV_X1 p9_mult_21_U822 ( .A(B3[11]), .ZN(p9_mult_21_n897) );
  INV_X1 p9_mult_21_U894 ( .A(B3[12]), .ZN(p9_mult_21_n879) );
  INV_X1 p9_mult_21_U453 ( .A(p9_mult_21_n901), .ZN(p9_mult_21_n899) );
  INV_X1 p9_mult_21_U859 ( .A(B3[9]), .ZN(p9_mult_21_n935) );
  INV_X1 p9_mult_21_U827 ( .A(p9_mult_21_n1092), .ZN(p9_mult_21_n863) );
  INV_X1 p9_mult_21_U863 ( .A(B3[10]), .ZN(p9_mult_21_n921) );
  INV_X1 p9_mult_21_U568 ( .A(p9_mult_21_n1063), .ZN(p9_mult_21_n862) );
  INV_X1 p9_mult_21_U816 ( .A(B3[13]), .ZN(p9_mult_21_n868) );
  INV_X1 p9_mult_21_U766 ( .A(p9_mult_21_n937), .ZN(p9_mult_21_n918) );
  INV_X1 p9_mult_21_U765 ( .A(p9_mult_21_n964), .ZN(p9_mult_21_n917) );
  OAI22_X1 p9_mult_21_U883 ( .A1(p9_mult_21_n1397), .A2(p9_mult_21_n987), .B1(
        reg4_reg[7]), .B2(reg4_reg[8]), .ZN(p9_mult_21_n964) );
  OAI22_X1 p9_mult_21_U874 ( .A1(p9_mult_21_n939), .A2(p9_mult_21_n1395), .B1(
        reg4_reg[10]), .B2(reg4_reg[9]), .ZN(p9_mult_21_n911) );
  XOR2_X1 p9_mult_21_U921 ( .A(p9_mult_21_n979), .B(p9_mult_21_n1003), .Z(
        p9_mult_21_n976) );
  XNOR2_X1 p9_mult_21_U645 ( .A(p9_mult_21_n1143), .B(p9_mult_21_n1177), .ZN(
        temp4[0]) );
  XNOR2_X1 p9_mult_21_U618 ( .A(p9_mult_21_n1140), .B(p9_mult_21_n1138), .ZN(
        temp4[1]) );
  XNOR2_X1 p9_mult_21_U620 ( .A(p9_mult_21_n1137), .B(p9_mult_21_n1139), .ZN(
        p9_mult_21_n1140) );
  XNOR2_X1 p9_mult_21_U592 ( .A(p9_mult_21_n1100), .B(p9_mult_21_n1104), .ZN(
        temp4[2]) );
  XNOR2_X1 p9_mult_21_U570 ( .A(p9_mult_21_n1067), .B(p9_mult_21_n1035), .ZN(
        temp4[3]) );
  XNOR2_X1 p9_mult_21_U589 ( .A(p9_mult_21_n1033), .B(p9_mult_21_n1034), .ZN(
        p9_mult_21_n1067) );
  XNOR2_X1 p9_mult_21_U543 ( .A(p9_mult_21_n1028), .B(p9_mult_21_n1032), .ZN(
        temp4[4]) );
  XNOR2_X1 p9_mult_21_U523 ( .A(p9_mult_21_n1002), .B(p9_mult_21_n976), .ZN(
        temp4[5]) );
  XNOR2_X1 p9_mult_21_U501 ( .A(p9_mult_21_n969), .B(p9_mult_21_n973), .ZN(
        temp4[6]) );
  XNOR2_X1 p9_mult_21_U485 ( .A(p9_mult_21_n948), .B(p9_mult_21_n928), .ZN(
        temp4[7]) );
  XNOR2_X1 p9_mult_21_U459 ( .A(p9_mult_21_n889), .B(p9_mult_21_n890), .ZN(
        p9_mult_21_n906) );
  XNOR2_X1 p9_mult_21_U469 ( .A(p9_mult_21_n909), .B(p9_mult_21_n925), .ZN(
        temp4[8]) );
  XNOR2_X1 p9_mult_21_U447 ( .A(p9_mult_21_n885), .B(p9_mult_21_n888), .ZN(
        temp4[10]) );
  XNOR2_X1 p9_mult_21_U439 ( .A(p9_mult_21_n876), .B(p9_mult_21_n871), .ZN(
        temp4[11]) );
  XNOR2_X1 p9_mult_21_U432 ( .A(p9_mult_21_n865), .B(p9_mult_21_n860), .ZN(
        temp4[12]) );
  AOI222_X1 p9_mult_21_U437 ( .A1(p9_mult_21_n872), .A2(p9_mult_21_n873), .B1(
        p9_mult_21_n872), .B2(p9_mult_21_n874), .C1(p9_mult_21_n873), .C2(
        p9_mult_21_n874), .ZN(p9_mult_21_n857) );
  AOI22_X1 p9_mult_21_U433 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n864), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n866), .ZN(p9_mult_21_n860) );
  AOI22_X1 p9_mult_21_U434 ( .A1(B3[13]), .A2(reg4_reg[13]), .B1(
        p9_mult_21_n867), .B2(p9_mult_21_n868), .ZN(p9_mult_21_n864) );
  XNOR2_X1 p9_mult_21_U440 ( .A(p9_mult_21_n874), .B(p9_mult_21_n875), .ZN(
        p9_mult_21_n877) );
  AOI22_X1 p9_mult_21_U441 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n866), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n878), .ZN(p9_mult_21_n875) );
  OAI22_X1 p9_mult_21_U442 ( .A1(p9_mult_21_n867), .A2(B3[12]), .B1(
        p9_mult_21_n879), .B2(reg4_reg[13]), .ZN(p9_mult_21_n866) );
  OAI21_X1 p9_mult_21_U443 ( .B1(p9_mult_21_n880), .B2(p9_mult_21_n881), .A(
        p9_mult_21_n882), .ZN(p9_mult_21_n872) );
  AOI222_X1 p9_mult_21_U449 ( .A1(p9_mult_21_n892), .A2(p9_mult_21_n893), .B1(
        p9_mult_21_n892), .B2(p9_mult_21_n894), .C1(p9_mult_21_n893), .C2(
        p9_mult_21_n894), .ZN(p9_mult_21_n883) );
  AOI222_X1 p9_mult_21_U468 ( .A1(p9_mult_21_n922), .A2(p9_mult_21_n923), .B1(
        p9_mult_21_n922), .B2(p9_mult_21_n924), .C1(p9_mult_21_n923), .C2(
        p9_mult_21_n924), .ZN(p9_mult_21_n889) );
  OAI22_X1 p9_mult_21_U460 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n902), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n912), .ZN(p9_mult_21_n893) );
  AOI222_X1 p9_mult_21_U462 ( .A1(p9_mult_21_n913), .A2(p9_mult_21_n914), .B1(
        p9_mult_21_n913), .B2(p9_mult_21_n900), .C1(p9_mult_21_n914), .C2(
        p9_mult_21_n900), .ZN(p9_mult_21_n892) );
  XNOR2_X1 p9_mult_21_U465 ( .A(p9_mult_21_n900), .B(p9_mult_21_n901), .ZN(
        p9_mult_21_n916) );
  XNOR2_X1 p9_mult_21_U472 ( .A(p9_mult_21_n932), .B(p9_mult_21_n924), .ZN(
        p9_mult_21_n909) );
  XNOR2_X1 p9_mult_21_U473 ( .A(p9_mult_21_n915), .B(p9_mult_21_n933), .ZN(
        p9_mult_21_n924) );
  AOI22_X1 p9_mult_21_U474 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n920), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n934), .ZN(p9_mult_21_n913) );
  OAI22_X1 p9_mult_21_U479 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n912), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n940), .ZN(p9_mult_21_n915) );
  OAI22_X1 p9_mult_21_U480 ( .A1(p9_mult_21_n905), .A2(p9_mult_21_n897), .B1(
        B3[11]), .B2(reg4_reg[11]), .ZN(p9_mult_21_n912) );
  XNOR2_X1 p9_mult_21_U481 ( .A(p9_mult_21_n922), .B(p9_mult_21_n923), .ZN(
        p9_mult_21_n932) );
  AOI222_X1 p9_mult_21_U482 ( .A1(p9_mult_21_n941), .A2(p9_mult_21_n942), .B1(
        p9_mult_21_n941), .B2(p9_mult_21_n943), .C1(p9_mult_21_n942), .C2(
        p9_mult_21_n943), .ZN(p9_mult_21_n923) );
  AOI222_X1 p9_mult_21_U483 ( .A1(p9_mult_21_n944), .A2(p9_mult_21_n945), .B1(
        p9_mult_21_n944), .B2(p9_mult_21_n946), .C1(p9_mult_21_n945), .C2(
        p9_mult_21_n946), .ZN(p9_mult_21_n922) );
  OAI21_X1 p9_mult_21_U486 ( .B1(p9_mult_21_n951), .B2(p9_mult_21_n952), .A(
        p9_mult_21_n953), .ZN(p9_mult_21_n944) );
  XNOR2_X1 p9_mult_21_U487 ( .A(p9_mult_21_n946), .B(p9_mult_21_n947), .ZN(
        p9_mult_21_n950) );
  AOI22_X1 p9_mult_21_U488 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n934), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n954), .ZN(p9_mult_21_n947) );
  AOI22_X1 p9_mult_21_U489 ( .A1(reg4_reg[13]), .A2(B3[8]), .B1(
        p9_mult_21_n955), .B2(p9_mult_21_n867), .ZN(p9_mult_21_n934) );
  AOI222_X1 p9_mult_21_U490 ( .A1(p9_mult_21_n956), .A2(p9_mult_21_n957), .B1(
        p9_mult_21_n956), .B2(p9_mult_21_n958), .C1(p9_mult_21_n957), .C2(
        p9_mult_21_n958), .ZN(p9_mult_21_n929) );
  OAI22_X1 p9_mult_21_U491 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n940), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n960), .ZN(p9_mult_21_n942) );
  OAI22_X1 p9_mult_21_U492 ( .A1(p9_mult_21_n905), .A2(p9_mult_21_n921), .B1(
        B3[10]), .B2(reg4_reg[11]), .ZN(p9_mult_21_n940) );
  AOI222_X1 p9_mult_21_U493 ( .A1(p9_mult_21_n961), .A2(p9_mult_21_n962), .B1(
        p9_mult_21_n961), .B2(p9_mult_21_n946), .C1(p9_mult_21_n962), .C2(
        p9_mult_21_n946), .ZN(p9_mult_21_n941) );
  OAI22_X1 p9_mult_21_U495 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n936), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n965), .ZN(p9_mult_21_n943) );
  AOI222_X1 p9_mult_21_U503 ( .A1(p9_mult_21_n977), .A2(p9_mult_21_n978), .B1(
        p9_mult_21_n977), .B2(p9_mult_21_n979), .C1(p9_mult_21_n978), .C2(
        p9_mult_21_n979), .ZN(p9_mult_21_n967) );
  XNOR2_X1 p9_mult_21_U504 ( .A(p9_mult_21_n980), .B(p9_mult_21_n972), .ZN(
        p9_mult_21_n969) );
  XNOR2_X1 p9_mult_21_U513 ( .A(p9_mult_21_n970), .B(p9_mult_21_n971), .ZN(
        p9_mult_21_n980) );
  AOI222_X1 p9_mult_21_U524 ( .A1(p9_mult_21_n1004), .A2(p9_mult_21_n1005), 
        .B1(p9_mult_21_n1004), .B2(p9_mult_21_n1006), .C1(p9_mult_21_n1005), 
        .C2(p9_mult_21_n1006), .ZN(p9_mult_21_n978) );
  AOI222_X1 p9_mult_21_U525 ( .A1(p9_mult_21_n1007), .A2(p9_mult_21_n1008), 
        .B1(p9_mult_21_n1007), .B2(p9_mult_21_n1009), .C1(p9_mult_21_n1008), 
        .C2(p9_mult_21_n1009), .ZN(p9_mult_21_n977) );
  AOI222_X1 p9_mult_21_U621 ( .A1(p9_mult_21_n1144), .A2(p9_mult_21_n1145), 
        .B1(p9_mult_21_n1144), .B2(p9_mult_21_n1146), .C1(p9_mult_21_n1145), 
        .C2(p9_mult_21_n1146), .ZN(p9_mult_21_n1139) );
  XNOR2_X1 p9_mult_21_U782 ( .A(p9_mult_21_n1359), .B(p9_mult_21_n1159), .ZN(
        p9_mult_21_n1145) );
  XNOR2_X1 p9_mult_21_U796 ( .A(p9_mult_21_n1160), .B(p9_mult_21_n1161), .ZN(
        p9_mult_21_n1359) );
  XNOR2_X1 p9_mult_21_U823 ( .A(p9_mult_21_n1377), .B(p9_mult_21_n1170), .ZN(
        p9_mult_21_n1146) );
  XNOR2_X1 p9_mult_21_U832 ( .A(p9_mult_21_n1169), .B(p9_mult_21_n1168), .ZN(
        p9_mult_21_n1377) );
  AOI222_X1 p9_mult_21_U836 ( .A1(p9_mult_21_n1351), .A2(p9_mult_21_n1353), 
        .B1(p9_mult_21_n1351), .B2(p9_mult_21_n1387), .C1(p9_mult_21_n1353), 
        .C2(p9_mult_21_n1387), .ZN(p9_mult_21_n1144) );
  AOI222_X1 p9_mult_21_U767 ( .A1(p9_mult_21_n1183), .A2(p9_mult_21_n1184), 
        .B1(p9_mult_21_n1183), .B2(p9_mult_21_n1182), .C1(p9_mult_21_n1184), 
        .C2(p9_mult_21_n1182), .ZN(p9_mult_21_n1142) );
  AOI222_X1 p9_mult_21_U768 ( .A1(p9_mult_21_n1324), .A2(p9_mult_21_n1325), 
        .B1(p9_mult_21_n1324), .B2(p9_mult_21_n1323), .C1(p9_mult_21_n1325), 
        .C2(p9_mult_21_n1323), .ZN(p9_mult_21_n1182) );
  XNOR2_X1 p9_mult_21_U648 ( .A(p9_mult_21_n1183), .B(p9_mult_21_n1184), .ZN(
        p9_mult_21_n1181) );
  XNOR2_X1 p9_mult_21_U781 ( .A(p9_mult_21_n1350), .B(p9_mult_21_n1351), .ZN(
        p9_mult_21_n1184) );
  XNOR2_X1 p9_mult_21_U847 ( .A(p9_mult_21_n1392), .B(p9_mult_21_n1385), .ZN(
        p9_mult_21_n1353) );
  AOI222_X1 p9_mult_21_U838 ( .A1(p9_mult_21_n1327), .A2(p9_mult_21_n1329), 
        .B1(p9_mult_21_n1327), .B2(p9_mult_21_n1328), .C1(p9_mult_21_n1329), 
        .C2(p9_mult_21_n1328), .ZN(p9_mult_21_n1352) );
  XNOR2_X1 p9_mult_21_U746 ( .A(p9_mult_21_n1322), .B(p9_mult_21_n1323), .ZN(
        p9_mult_21_n1186) );
  XNOR2_X1 p9_mult_21_U769 ( .A(p9_mult_21_n1343), .B(p9_mult_21_n1344), .ZN(
        p9_mult_21_n1341) );
  XNOR2_X1 p9_mult_21_U747 ( .A(p9_mult_21_n1324), .B(p9_mult_21_n1325), .ZN(
        p9_mult_21_n1322) );
  AOI222_X1 p9_mult_21_U770 ( .A1(p9_mult_21_n1337), .A2(p9_mult_21_n1336), 
        .B1(p9_mult_21_n1337), .B2(p9_mult_21_n1335), .C1(p9_mult_21_n1336), 
        .C2(p9_mult_21_n1335), .ZN(p9_mult_21_n1325) );
  AOI222_X1 p9_mult_21_U774 ( .A1(p9_mult_21_n1205), .A2(p9_mult_21_n1206), 
        .B1(p9_mult_21_n1205), .B2(p9_mult_21_n1204), .C1(p9_mult_21_n1206), 
        .C2(p9_mult_21_n1204), .ZN(p9_mult_21_n1324) );
  XNOR2_X1 p9_mult_21_U748 ( .A(p9_mult_21_n1328), .B(p9_mult_21_n1329), .ZN(
        p9_mult_21_n1326) );
  AOI222_X1 p9_mult_21_U749 ( .A1(p9_mult_21_n1199), .A2(p9_mult_21_n1202), 
        .B1(p9_mult_21_n1199), .B2(p9_mult_21_n1201), .C1(p9_mult_21_n1202), 
        .C2(p9_mult_21_n1201), .ZN(p9_mult_21_n1185) );
  AOI222_X1 p9_mult_21_U651 ( .A1(p9_mult_21_n1191), .A2(p9_mult_21_n1192), 
        .B1(p9_mult_21_n1191), .B2(p9_mult_21_n1193), .C1(p9_mult_21_n1192), 
        .C2(p9_mult_21_n1193), .ZN(p9_mult_21_n1190) );
  XNOR2_X1 p9_mult_21_U654 ( .A(p9_mult_21_n1198), .B(p9_mult_21_n1193), .ZN(
        p9_mult_21_n1197) );
  XNOR2_X1 p9_mult_21_U758 ( .A(p9_mult_21_n1334), .B(p9_mult_21_n1335), .ZN(
        p9_mult_21_n1202) );
  XNOR2_X1 p9_mult_21_U759 ( .A(p9_mult_21_n1336), .B(p9_mult_21_n1337), .ZN(
        p9_mult_21_n1334) );
  OAI22_X1 p9_mult_21_U840 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n1094), .B1(
        B3[4]), .B2(reg4_reg[7]), .ZN(p9_mult_21_n1346) );
  OAI222_X1 p9_mult_21_U751 ( .A1(p9_mult_21_n1314), .A2(p9_mult_21_n1315), 
        .B1(p9_mult_21_n1314), .B2(p9_mult_21_n1313), .C1(p9_mult_21_n1315), 
        .C2(p9_mult_21_n1313), .ZN(p9_mult_21_n1330) );
  NOR2_X1 p9_mult_21_U760 ( .A1(p9_mult_21_n1308), .A2(p9_mult_21_n1307), .ZN(
        p9_mult_21_n1199) );
  XNOR2_X1 p9_mult_21_U655 ( .A(p9_mult_21_n1203), .B(p9_mult_21_n1204), .ZN(
        p9_mult_21_n1192) );
  XNOR2_X1 p9_mult_21_U656 ( .A(p9_mult_21_n1205), .B(p9_mult_21_n1206), .ZN(
        p9_mult_21_n1203) );
  OAI22_X1 p9_mult_21_U779 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1349), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1340), .ZN(p9_mult_21_n1205) );
  AOI222_X1 p9_mult_21_U657 ( .A1(p9_mult_21_n1207), .A2(p9_mult_21_n1208), 
        .B1(p9_mult_21_n1207), .B2(p9_mult_21_n1209), .C1(p9_mult_21_n1208), 
        .C2(p9_mult_21_n1209), .ZN(p9_mult_21_n1194) );
  AOI222_X1 p9_mult_21_U658 ( .A1(p9_mult_21_n1210), .A2(p9_mult_21_n1211), 
        .B1(p9_mult_21_n1210), .B2(p9_mult_21_n1212), .C1(p9_mult_21_n1211), 
        .C2(p9_mult_21_n1212), .ZN(p9_mult_21_n1196) );
  XNOR2_X1 p9_mult_21_U663 ( .A(p9_mult_21_n1224), .B(p9_mult_21_n1225), .ZN(
        p9_mult_21_n1217) );
  XNOR2_X1 p9_mult_21_U664 ( .A(p9_mult_21_n1226), .B(p9_mult_21_n1227), .ZN(
        p9_mult_21_n1224) );
  XNOR2_X1 p9_mult_21_U665 ( .A(p9_mult_21_n1219), .B(p9_mult_21_n1216), .ZN(
        p9_mult_21_n1223) );
  AOI222_X1 p9_mult_21_U666 ( .A1(p9_mult_21_n1232), .A2(p9_mult_21_n1233), 
        .B1(p9_mult_21_n1232), .B2(p9_mult_21_n1234), .C1(p9_mult_21_n1233), 
        .C2(p9_mult_21_n1234), .ZN(p9_mult_21_n1219) );
  XNOR2_X1 p9_mult_21_U670 ( .A(p9_mult_21_n1232), .B(p9_mult_21_n1234), .ZN(
        p9_mult_21_n1242) );
  XNOR2_X1 p9_mult_21_U673 ( .A(p9_mult_21_n1250), .B(p9_mult_21_n1251), .ZN(
        p9_mult_21_n1237) );
  AOI222_X1 p9_mult_21_U674 ( .A1(p9_mult_21_n1252), .A2(p9_mult_21_n1253), 
        .B1(p9_mult_21_n1252), .B2(p9_mult_21_n1254), .C1(p9_mult_21_n1253), 
        .C2(p9_mult_21_n1254), .ZN(p9_mult_21_n1235) );
  XNOR2_X1 p9_mult_21_U716 ( .A(p9_mult_21_n1302), .B(p9_mult_21_n1254), .ZN(
        p9_mult_21_n1258) );
  NOR2_X1 p9_mult_21_U417 ( .A1(B3[5]), .A2(p9_mult_21_n1245), .ZN(
        p9_mult_21_n844) );
  XNOR2_X1 p9_mult_21_U718 ( .A(p9_mult_21_n1253), .B(p9_mult_21_n1252), .ZN(
        p9_mult_21_n1302) );
  NOR2_X1 p9_mult_21_U411 ( .A1(B3[4]), .A2(p9_mult_21_n1245), .ZN(
        p9_mult_21_n838) );
  OAI22_X1 p9_mult_21_U697 ( .A1(B3[1]), .A2(p9_mult_21_n1294), .B1(
        p9_mult_21_n1295), .B2(p9_mult_21_n1244), .ZN(p9_mult_21_n1293) );
  NOR2_X1 p9_mult_21_U415 ( .A1(B3[2]), .A2(p9_mult_21_n1245), .ZN(
        p9_mult_21_n842) );
  NOR2_X1 p9_mult_21_U413 ( .A1(B3[3]), .A2(p9_mult_21_n1245), .ZN(
        p9_mult_21_n840) );
  XNOR2_X1 p9_mult_21_U724 ( .A(p9_mult_21_n1305), .B(p9_mult_21_n1208), .ZN(
        p9_mult_21_n1212) );
  AOI21_X1 p9_mult_21_U761 ( .B1(p9_mult_21_n1338), .B2(p9_mult_21_n917), .A(
        p9_mult_21_n1339), .ZN(p9_mult_21_n1307) );
  AOI222_X1 p9_mult_21_U727 ( .A1(p9_mult_21_n1227), .A2(p9_mult_21_n1226), 
        .B1(p9_mult_21_n1227), .B2(p9_mult_21_n1225), .C1(p9_mult_21_n1226), 
        .C2(p9_mult_21_n1225), .ZN(p9_mult_21_n1309) );
  XNOR2_X1 p9_mult_21_U732 ( .A(p9_mult_21_n1211), .B(p9_mult_21_n1210), .ZN(
        p9_mult_21_n1304) );
  XNOR2_X1 p9_mult_21_U733 ( .A(p9_mult_21_n1314), .B(p9_mult_21_n1315), .ZN(
        p9_mult_21_n1312) );
  AOI222_X1 p9_mult_21_U734 ( .A1(p9_mult_21_n1231), .A2(p9_mult_21_n1230), 
        .B1(p9_mult_21_n1231), .B2(p9_mult_21_n1228), .C1(p9_mult_21_n1230), 
        .C2(p9_mult_21_n1228), .ZN(p9_mult_21_n1211) );
  OAI22_X1 p9_mult_21_U757 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n1175), .B1(
        B3[2]), .B2(reg4_reg[7]), .ZN(p9_mult_21_n1317) );
  NOR2_X1 p9_mult_21_U738 ( .A1(p9_mult_21_n1251), .A2(p9_mult_21_n1250), .ZN(
        p9_mult_21_n1231) );
  XNOR2_X1 p9_mult_21_U593 ( .A(p9_mult_21_n1105), .B(p9_mult_21_n1103), .ZN(
        p9_mult_21_n1099) );
  XNOR2_X1 p9_mult_21_U609 ( .A(p9_mult_21_n1101), .B(p9_mult_21_n1102), .ZN(
        p9_mult_21_n1105) );
  AOI222_X1 p9_mult_21_U616 ( .A1(p9_mult_21_n1134), .A2(p9_mult_21_n1135), 
        .B1(p9_mult_21_n1134), .B2(p9_mult_21_n1136), .C1(p9_mult_21_n1135), 
        .C2(p9_mult_21_n1136), .ZN(p9_mult_21_n1098) );
  AOI222_X1 p9_mult_21_U631 ( .A1(p9_mult_21_n1159), .A2(p9_mult_21_n1160), 
        .B1(p9_mult_21_n1159), .B2(p9_mult_21_n1161), .C1(p9_mult_21_n1160), 
        .C2(p9_mult_21_n1161), .ZN(p9_mult_21_n1136) );
  XNOR2_X1 p9_mult_21_U799 ( .A(p9_mult_21_n1155), .B(p9_mult_21_n1156), .ZN(
        p9_mult_21_n1367) );
  XNOR2_X1 p9_mult_21_U811 ( .A(p9_mult_21_n1154), .B(p9_mult_21_n1372), .ZN(
        p9_mult_21_n1160) );
  AOI222_X1 p9_mult_21_U783 ( .A1(p9_mult_21_n1357), .A2(p9_mult_21_n1356), 
        .B1(p9_mult_21_n1357), .B2(p9_mult_21_n1354), .C1(p9_mult_21_n1356), 
        .C2(p9_mult_21_n1354), .ZN(p9_mult_21_n1159) );
  OAI222_X1 p9_mult_21_U786 ( .A1(p9_mult_21_n1343), .A2(p9_mult_21_n1344), 
        .B1(p9_mult_21_n1343), .B2(p9_mult_21_n1342), .C1(p9_mult_21_n1344), 
        .C2(p9_mult_21_n1342), .ZN(p9_mult_21_n1362) );
  OAI22_X1 p9_mult_21_U787 ( .A1(p9_mult_21_n1244), .A2(p9_mult_21_n1363), 
        .B1(p9_mult_21_n1294), .B2(p9_mult_21_n1345), .ZN(p9_mult_21_n1342) );
  OAI22_X1 p9_mult_21_U793 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1364), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1349), .ZN(p9_mult_21_n1343) );
  OAI22_X1 p9_mult_21_U794 ( .A1(p9_mult_21_n939), .A2(p9_mult_21_n1175), .B1(
        B3[2]), .B2(reg4_reg[9]), .ZN(p9_mult_21_n1349) );
  NOR2_X1 p9_mult_21_U795 ( .A1(p9_mult_21_n1365), .A2(p9_mult_21_n1366), .ZN(
        p9_mult_21_n1357) );
  AOI21_X1 p9_mult_21_U845 ( .B1(p9_mult_21_n1390), .B2(p9_mult_21_n880), .A(
        p9_mult_21_n1391), .ZN(p9_mult_21_n1366) );
  XNOR2_X1 p9_mult_21_U632 ( .A(p9_mult_21_n1162), .B(p9_mult_21_n1133), .ZN(
        p9_mult_21_n1134) );
  XNOR2_X1 p9_mult_21_U638 ( .A(p9_mult_21_n1131), .B(p9_mult_21_n1132), .ZN(
        p9_mult_21_n1162) );
  AOI222_X1 p9_mult_21_U591 ( .A1(p9_mult_21_n1101), .A2(p9_mult_21_n1102), 
        .B1(p9_mult_21_n1101), .B2(p9_mult_21_n1103), .C1(p9_mult_21_n1102), 
        .C2(p9_mult_21_n1103), .ZN(p9_mult_21_n1033) );
  XNOR2_X1 p9_mult_21_U610 ( .A(p9_mult_21_n1122), .B(p9_mult_21_n1097), .ZN(
        p9_mult_21_n1102) );
  XNOR2_X1 p9_mult_21_U612 ( .A(p9_mult_21_n1095), .B(p9_mult_21_n1096), .ZN(
        p9_mult_21_n1122) );
  AOI222_X1 p9_mult_21_U615 ( .A1(p9_mult_21_n1131), .A2(p9_mult_21_n1132), 
        .B1(p9_mult_21_n1131), .B2(p9_mult_21_n1133), .C1(p9_mult_21_n1132), 
        .C2(p9_mult_21_n1133), .ZN(p9_mult_21_n1101) );
  AOI222_X1 p9_mult_21_U639 ( .A1(p9_mult_21_n1168), .A2(p9_mult_21_n1169), 
        .B1(p9_mult_21_n1168), .B2(p9_mult_21_n1170), .C1(p9_mult_21_n1169), 
        .C2(p9_mult_21_n1170), .ZN(p9_mult_21_n1132) );
  XNOR2_X1 p9_mult_21_U824 ( .A(p9_mult_21_n1172), .B(p9_mult_21_n1173), .ZN(
        p9_mult_21_n1170) );
  AOI222_X1 p9_mult_21_U834 ( .A1(p9_mult_21_n1383), .A2(p9_mult_21_n1384), 
        .B1(p9_mult_21_n1383), .B2(p9_mult_21_n1385), .C1(p9_mult_21_n1384), 
        .C2(p9_mult_21_n1385), .ZN(p9_mult_21_n1169) );
  AOI22_X1 p9_mult_21_U849 ( .A1(reg4_reg[7]), .A2(p9_mult_21_n1062), .B1(
        B3[5]), .B2(p9_mult_21_n987), .ZN(p9_mult_21_n1388) );
  AOI22_X1 p9_mult_21_U866 ( .A1(p9_mult_21_n880), .A2(p9_mult_21_n1371), .B1(
        p9_mult_21_n881), .B2(p9_mult_21_n1390), .ZN(p9_mult_21_n1386) );
  AOI222_X1 p9_mult_21_U833 ( .A1(p9_mult_21_n1380), .A2(p9_mult_21_n1381), 
        .B1(p9_mult_21_n1380), .B2(p9_mult_21_n1382), .C1(p9_mult_21_n1381), 
        .C2(p9_mult_21_n1382), .ZN(p9_mult_21_n1168) );
  OAI22_X1 p9_mult_21_U876 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1368), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1364), .ZN(p9_mult_21_n1381) );
  AOI222_X1 p9_mult_21_U545 ( .A1(p9_mult_21_n1036), .A2(p9_mult_21_n1037), 
        .B1(p9_mult_21_n1036), .B2(p9_mult_21_n1038), .C1(p9_mult_21_n1037), 
        .C2(p9_mult_21_n1038), .ZN(p9_mult_21_n1026) );
  AOI222_X1 p9_mult_21_U576 ( .A1(p9_mult_21_n1077), .A2(p9_mult_21_n1078), 
        .B1(p9_mult_21_n1077), .B2(p9_mult_21_n1079), .C1(p9_mult_21_n1078), 
        .C2(p9_mult_21_n1079), .ZN(p9_mult_21_n1036) );
  XNOR2_X1 p9_mult_21_U604 ( .A(p9_mult_21_n1071), .B(p9_mult_21_n1072), .ZN(
        p9_mult_21_n1117) );
  AOI222_X1 p9_mult_21_U594 ( .A1(p9_mult_21_n1107), .A2(p9_mult_21_n1108), 
        .B1(p9_mult_21_n1107), .B2(p9_mult_21_n1109), .C1(p9_mult_21_n1108), 
        .C2(p9_mult_21_n1109), .ZN(p9_mult_21_n1077) );
  XNOR2_X1 p9_mult_21_U622 ( .A(p9_mult_21_n1123), .B(p9_mult_21_n1124), .ZN(
        p9_mult_21_n1109) );
  AOI222_X1 p9_mult_21_U629 ( .A1(p9_mult_21_n1155), .A2(p9_mult_21_n1156), 
        .B1(p9_mult_21_n1155), .B2(p9_mult_21_n1157), .C1(p9_mult_21_n1156), 
        .C2(p9_mult_21_n1157), .ZN(p9_mult_21_n1108) );
  OAI22_X1 p9_mult_21_U797 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1164), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1368), .ZN(p9_mult_21_n1158) );
  OAI22_X1 p9_mult_21_U880 ( .A1(p9_mult_21_n939), .A2(p9_mult_21_n1094), .B1(
        B3[4]), .B2(reg4_reg[9]), .ZN(p9_mult_21_n1368) );
  AOI22_X1 p9_mult_21_U800 ( .A1(p9_mult_21_n1021), .A2(p9_mult_21_n1150), 
        .B1(p9_mult_21_n1022), .B2(p9_mult_21_n1369), .ZN(p9_mult_21_n1156) );
  AOI22_X1 p9_mult_21_U809 ( .A1(p9_mult_21_n880), .A2(p9_mult_21_n1149), .B1(
        p9_mult_21_n881), .B2(p9_mult_21_n1371), .ZN(p9_mult_21_n1155) );
  AOI22_X1 p9_mult_21_U871 ( .A1(reg4_reg[11]), .A2(B3[2]), .B1(
        p9_mult_21_n1175), .B2(p9_mult_21_n905), .ZN(p9_mult_21_n1371) );
  OAI222_X1 p9_mult_21_U628 ( .A1(p9_mult_21_n1152), .A2(p9_mult_21_n1153), 
        .B1(p9_mult_21_n1152), .B2(p9_mult_21_n1154), .C1(p9_mult_21_n1153), 
        .C2(p9_mult_21_n1154), .ZN(p9_mult_21_n1151) );
  OAI22_X1 p9_mult_21_U852 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n1025), .B1(
        B3[6]), .B2(reg4_reg[7]), .ZN(p9_mult_21_n1375) );
  OAI22_X1 p9_mult_21_U812 ( .A1(p9_mult_21_n1244), .A2(p9_mult_21_n1373), 
        .B1(p9_mult_21_n1294), .B2(p9_mult_21_n1374), .ZN(p9_mult_21_n1152) );
  XNOR2_X1 p9_mult_21_U546 ( .A(p9_mult_21_n1040), .B(p9_mult_21_n1006), .ZN(
        p9_mult_21_n1031) );
  XNOR2_X1 p9_mult_21_U547 ( .A(p9_mult_21_n1018), .B(p9_mult_21_n1041), .ZN(
        p9_mult_21_n1006) );
  XNOR2_X1 p9_mult_21_U548 ( .A(p9_mult_21_n993), .B(p9_mult_21_n1017), .ZN(
        p9_mult_21_n1041) );
  XNOR2_X1 p9_mult_21_U556 ( .A(p9_mult_21_n1004), .B(p9_mult_21_n1005), .ZN(
        p9_mult_21_n1040) );
  AOI222_X1 p9_mult_21_U557 ( .A1(p9_mult_21_n1048), .A2(p9_mult_21_n1049), 
        .B1(p9_mult_21_n1048), .B2(p9_mult_21_n1050), .C1(p9_mult_21_n1049), 
        .C2(p9_mult_21_n1050), .ZN(p9_mult_21_n1005) );
  AOI222_X1 p9_mult_21_U558 ( .A1(p9_mult_21_n1051), .A2(p9_mult_21_n1052), 
        .B1(p9_mult_21_n1051), .B2(p9_mult_21_n1053), .C1(p9_mult_21_n1052), 
        .C2(p9_mult_21_n1053), .ZN(p9_mult_21_n1004) );
  OAI222_X1 p9_mult_21_U572 ( .A1(p9_mult_21_n1071), .A2(p9_mult_21_n1072), 
        .B1(p9_mult_21_n1071), .B2(p9_mult_21_n1073), .C1(p9_mult_21_n1072), 
        .C2(p9_mult_21_n1073), .ZN(p9_mult_21_n1070) );
  OAI22_X1 p9_mult_21_U602 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1087), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1118), .ZN(p9_mult_21_n1073) );
  OAI22_X1 p9_mult_21_U606 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n935), .B1(
        B3[9]), .B2(reg4_reg[7]), .ZN(p9_mult_21_n1076) );
  OAI22_X1 p9_mult_21_U607 ( .A1(p9_mult_21_n1063), .A2(p9_mult_21_n1093), 
        .B1(p9_mult_21_n1092), .B2(p9_mult_21_n1120), .ZN(p9_mult_21_n1071) );
  AOI222_X1 p9_mult_21_U573 ( .A1(p9_mult_21_n1074), .A2(p9_mult_21_n1075), 
        .B1(p9_mult_21_n1074), .B2(p9_mult_21_n1066), .C1(p9_mult_21_n1075), 
        .C2(p9_mult_21_n1066), .ZN(p9_mult_21_n1051) );
  AOI22_X1 p9_mult_21_U600 ( .A1(p9_mult_21_n880), .A2(p9_mult_21_n1086), .B1(
        p9_mult_21_n881), .B2(p9_mult_21_n1116), .ZN(p9_mult_21_n1075) );
  AOI22_X1 p9_mult_21_U595 ( .A1(p9_mult_21_n1021), .A2(p9_mult_21_n1084), 
        .B1(p9_mult_21_n1022), .B2(p9_mult_21_n1111), .ZN(p9_mult_21_n1074) );
  XNOR2_X1 p9_mult_21_U560 ( .A(p9_mult_21_n1057), .B(p9_mult_21_n1009), .ZN(
        p9_mult_21_n1030) );
  AOI22_X1 p9_mult_21_U561 ( .A1(p9_mult_21_n917), .A2(p9_mult_21_n1013), .B1(
        p9_mult_21_n918), .B2(p9_mult_21_n1058), .ZN(p9_mult_21_n1009) );
  XNOR2_X1 p9_mult_21_U564 ( .A(p9_mult_21_n1007), .B(p9_mult_21_n1008), .ZN(
        p9_mult_21_n1057) );
  AOI22_X1 p9_mult_21_U565 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n1024), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n1060), .ZN(p9_mult_21_n1008) );
  AOI222_X1 p9_mult_21_U569 ( .A1(p9_mult_21_n1064), .A2(p9_mult_21_n1065), 
        .B1(p9_mult_21_n1064), .B2(p9_mult_21_n1066), .C1(p9_mult_21_n1065), 
        .C2(p9_mult_21_n1066), .ZN(p9_mult_21_n1007) );
  AOI222_X1 p9_mult_21_U559 ( .A1(p9_mult_21_n1054), .A2(p9_mult_21_n1055), 
        .B1(p9_mult_21_n1054), .B2(p9_mult_21_n1056), .C1(p9_mult_21_n1055), 
        .C2(p9_mult_21_n1056), .ZN(p9_mult_21_n1029) );
  OAI22_X1 p9_mult_21_U580 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n1047), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n1085), .ZN(p9_mult_21_n1048) );
  AOI22_X1 p9_mult_21_U601 ( .A1(reg4_reg[11]), .A2(B3[5]), .B1(
        p9_mult_21_n1062), .B2(p9_mult_21_n905), .ZN(p9_mult_21_n1086) );
  OAI22_X1 p9_mult_21_U583 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1059), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1087), .ZN(p9_mult_21_n1050) );
  OAI22_X1 p9_mult_21_U603 ( .A1(p9_mult_21_n939), .A2(p9_mult_21_n983), .B1(
        B3[7]), .B2(reg4_reg[9]), .ZN(p9_mult_21_n1087) );
  OAI22_X1 p9_mult_21_U584 ( .A1(p9_mult_21_n939), .A2(p9_mult_21_n955), .B1(
        B3[8]), .B2(reg4_reg[9]), .ZN(p9_mult_21_n1059) );
  OAI22_X1 p9_mult_21_U586 ( .A1(p9_mult_21_n1063), .A2(p9_mult_21_n1061), 
        .B1(p9_mult_21_n1092), .B2(p9_mult_21_n1093), .ZN(p9_mult_21_n1065) );
  AOI22_X1 p9_mult_21_U587 ( .A1(reg4_reg[13]), .A2(p9_mult_21_n1094), .B1(
        B3[4]), .B2(p9_mult_21_n867), .ZN(p9_mult_21_n1061) );
  OAI21_X1 p9_mult_21_U597 ( .B1(p9_mult_21_n1112), .B2(p9_mult_21_n1113), .A(
        p9_mult_21_n1114), .ZN(p9_mult_21_n1066) );
  NAND2_X1 p9_mult_21_U598 ( .A1(p9_mult_21_n1089), .A2(p9_mult_21_n1091), 
        .ZN(p9_mult_21_n1114) );
  AOI222_X1 p9_mult_21_U588 ( .A1(p9_mult_21_n1095), .A2(p9_mult_21_n1096), 
        .B1(p9_mult_21_n1095), .B2(p9_mult_21_n1097), .C1(p9_mult_21_n1096), 
        .C2(p9_mult_21_n1097), .ZN(p9_mult_21_n1054) );
  AOI22_X1 p9_mult_21_U623 ( .A1(p9_mult_21_n880), .A2(p9_mult_21_n1116), .B1(
        p9_mult_21_n881), .B2(p9_mult_21_n1149), .ZN(p9_mult_21_n1124) );
  AOI22_X1 p9_mult_21_U624 ( .A1(reg4_reg[11]), .A2(B3[4]), .B1(
        p9_mult_21_n1094), .B2(p9_mult_21_n905), .ZN(p9_mult_21_n1116) );
  AOI22_X1 p9_mult_21_U625 ( .A1(p9_mult_21_n1021), .A2(p9_mult_21_n1111), 
        .B1(p9_mult_21_n1022), .B2(p9_mult_21_n1150), .ZN(p9_mult_21_n1123) );
  AOI222_X1 p9_mult_21_U613 ( .A1(p9_mult_21_n1125), .A2(p9_mult_21_n1126), 
        .B1(p9_mult_21_n1125), .B2(p9_mult_21_n1127), .C1(p9_mult_21_n1126), 
        .C2(p9_mult_21_n1127), .ZN(p9_mult_21_n1096) );
  OAI22_X1 p9_mult_21_U633 ( .A1(p9_mult_21_n964), .A2(p9_mult_21_n1118), .B1(
        p9_mult_21_n937), .B2(p9_mult_21_n1164), .ZN(p9_mult_21_n1126) );
  AOI22_X1 p9_mult_21_U798 ( .A1(reg4_reg[9]), .A2(p9_mult_21_n1062), .B1(
        B3[5]), .B2(p9_mult_21_n939), .ZN(p9_mult_21_n1164) );
  OAI22_X1 p9_mult_21_U634 ( .A1(p9_mult_21_n939), .A2(p9_mult_21_n1025), .B1(
        B3[6]), .B2(reg4_reg[9]), .ZN(p9_mult_21_n1118) );
  AOI222_X1 p9_mult_21_U614 ( .A1(p9_mult_21_n1128), .A2(p9_mult_21_n1129), 
        .B1(p9_mult_21_n1128), .B2(p9_mult_21_n1130), .C1(p9_mult_21_n1129), 
        .C2(p9_mult_21_n1130), .ZN(p9_mult_21_n1095) );
  AOI22_X1 p9_mult_21_U818 ( .A1(reg4_reg[7]), .A2(p9_mult_21_n983), .B1(B3[7]), .B2(p9_mult_21_n987), .ZN(p9_mult_21_n1176) );
  OAI22_X1 p9_mult_21_U644 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n955), .B1(
        B3[8]), .B2(reg4_reg[7]), .ZN(p9_mult_21_n1119) );
  OAI22_X1 p9_mult_21_U641 ( .A1(p9_mult_21_n1063), .A2(p9_mult_21_n1120), 
        .B1(p9_mult_21_n1092), .B2(p9_mult_21_n1174), .ZN(p9_mult_21_n1129) );
  OAI22_X1 p9_mult_21_U642 ( .A1(p9_mult_21_n867), .A2(p9_mult_21_n1175), .B1(
        B3[2]), .B2(reg4_reg[13]), .ZN(p9_mult_21_n1120) );
  OAI21_X1 p9_mult_21_U825 ( .B1(p9_mult_21_n1174), .B2(p9_mult_21_n1063), .A(
        p9_mult_21_n1378), .ZN(p9_mult_21_n1173) );
  AOI221_X1 p9_mult_21_U829 ( .B1(p9_mult_21_n1092), .B2(p9_mult_21_n1063), 
        .C1(p9_mult_21_n1092), .C2(B3[0]), .A(p9_mult_21_n867), .ZN(
        p9_mult_21_n1172) );
  AOI222_X1 p9_mult_21_U500 ( .A1(p9_mult_21_n970), .A2(p9_mult_21_n971), .B1(
        p9_mult_21_n970), .B2(p9_mult_21_n972), .C1(p9_mult_21_n971), .C2(
        p9_mult_21_n972), .ZN(p9_mult_21_n926) );
  XNOR2_X1 p9_mult_21_U505 ( .A(p9_mult_21_n963), .B(p9_mult_21_n981), .ZN(
        p9_mult_21_n972) );
  AOI22_X1 p9_mult_21_U506 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n954), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n982), .ZN(p9_mult_21_n961) );
  OAI22_X1 p9_mult_21_U507 ( .A1(p9_mult_21_n867), .A2(B3[7]), .B1(
        p9_mult_21_n983), .B2(reg4_reg[13]), .ZN(p9_mult_21_n954) );
  OAI21_X1 p9_mult_21_U508 ( .B1(p9_mult_21_n984), .B2(p9_mult_21_n985), .A(
        p9_mult_21_n986), .ZN(p9_mult_21_n946) );
  NAND2_X1 p9_mult_21_U509 ( .A1(p9_mult_21_n951), .A2(p9_mult_21_n953), .ZN(
        p9_mult_21_n986) );
  AOI22_X1 p9_mult_21_U510 ( .A1(B3[13]), .A2(reg4_reg[7]), .B1(
        p9_mult_21_n987), .B2(p9_mult_21_n868), .ZN(p9_mult_21_n953) );
  OAI22_X1 p9_mult_21_U511 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n960), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n988), .ZN(p9_mult_21_n963) );
  OAI22_X1 p9_mult_21_U512 ( .A1(p9_mult_21_n905), .A2(p9_mult_21_n935), .B1(
        B3[9]), .B2(reg4_reg[11]), .ZN(p9_mult_21_n960) );
  XNOR2_X1 p9_mult_21_U514 ( .A(p9_mult_21_n956), .B(p9_mult_21_n989), .ZN(
        p9_mult_21_n971) );
  XNOR2_X1 p9_mult_21_U515 ( .A(p9_mult_21_n957), .B(p9_mult_21_n958), .ZN(
        p9_mult_21_n989) );
  AOI22_X1 p9_mult_21_U516 ( .A1(p9_mult_21_n917), .A2(p9_mult_21_n966), .B1(
        p9_mult_21_n918), .B2(p9_mult_21_n990), .ZN(p9_mult_21_n958) );
  OAI22_X1 p9_mult_21_U517 ( .A1(p9_mult_21_n939), .A2(B3[11]), .B1(
        p9_mult_21_n897), .B2(reg4_reg[9]), .ZN(p9_mult_21_n966) );
  AOI222_X1 p9_mult_21_U518 ( .A1(p9_mult_21_n991), .A2(p9_mult_21_n992), .B1(
        p9_mult_21_n991), .B2(p9_mult_21_n993), .C1(p9_mult_21_n992), .C2(
        p9_mult_21_n993), .ZN(p9_mult_21_n957) );
  AOI222_X1 p9_mult_21_U520 ( .A1(p9_mult_21_n995), .A2(p9_mult_21_n996), .B1(
        p9_mult_21_n995), .B2(p9_mult_21_n997), .C1(p9_mult_21_n996), .C2(
        p9_mult_21_n997), .ZN(p9_mult_21_n956) );
  AOI222_X1 p9_mult_21_U522 ( .A1(p9_mult_21_n999), .A2(p9_mult_21_n1000), 
        .B1(p9_mult_21_n999), .B2(p9_mult_21_n1001), .C1(p9_mult_21_n1000), 
        .C2(p9_mult_21_n1001), .ZN(p9_mult_21_n970) );
  OAI21_X1 p9_mult_21_U536 ( .B1(p9_mult_21_n1021), .B2(p9_mult_21_n1022), .A(
        p9_mult_21_n1023), .ZN(p9_mult_21_n991) );
  XNOR2_X1 p9_mult_21_U537 ( .A(p9_mult_21_n993), .B(p9_mult_21_n994), .ZN(
        p9_mult_21_n1020) );
  AOI22_X1 p9_mult_21_U538 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n982), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n1024), .ZN(p9_mult_21_n994) );
  OAI22_X1 p9_mult_21_U567 ( .A1(p9_mult_21_n867), .A2(B3[5]), .B1(
        p9_mult_21_n1062), .B2(reg4_reg[13]), .ZN(p9_mult_21_n1024) );
  AOI22_X1 p9_mult_21_U539 ( .A1(reg4_reg[13]), .A2(B3[6]), .B1(
        p9_mult_21_n1025), .B2(p9_mult_21_n867), .ZN(p9_mult_21_n982) );
  XNOR2_X1 p9_mult_21_U526 ( .A(p9_mult_21_n998), .B(p9_mult_21_n996), .ZN(
        p9_mult_21_n1011) );
  OAI22_X1 p9_mult_21_U527 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n988), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n1012), .ZN(p9_mult_21_n996) );
  OAI22_X1 p9_mult_21_U528 ( .A1(p9_mult_21_n905), .A2(p9_mult_21_n955), .B1(
        B3[8]), .B2(reg4_reg[11]), .ZN(p9_mult_21_n988) );
  AOI22_X1 p9_mult_21_U529 ( .A1(p9_mult_21_n917), .A2(p9_mult_21_n990), .B1(
        p9_mult_21_n918), .B2(p9_mult_21_n1013), .ZN(p9_mult_21_n998) );
  OAI22_X1 p9_mult_21_U563 ( .A1(p9_mult_21_n939), .A2(B3[9]), .B1(
        p9_mult_21_n935), .B2(reg4_reg[9]), .ZN(p9_mult_21_n1013) );
  OAI22_X1 p9_mult_21_U530 ( .A1(p9_mult_21_n939), .A2(B3[10]), .B1(
        p9_mult_21_n921), .B2(reg4_reg[9]), .ZN(p9_mult_21_n990) );
  AOI22_X1 p9_mult_21_U532 ( .A1(B3[12]), .A2(p9_mult_21_n987), .B1(
        reg4_reg[7]), .B2(p9_mult_21_n879), .ZN(p9_mult_21_n984) );
  OAI222_X1 p9_mult_21_U534 ( .A1(p9_mult_21_n1017), .A2(p9_mult_21_n1018), 
        .B1(p9_mult_21_n1017), .B2(p9_mult_21_n1019), .C1(p9_mult_21_n1018), 
        .C2(p9_mult_21_n1019), .ZN(p9_mult_21_n1016) );
  OAI21_X1 p9_mult_21_U551 ( .B1(p9_mult_21_n1043), .B2(p9_mult_21_n1044), .A(
        p9_mult_21_n1045), .ZN(p9_mult_21_n993) );
  NAND2_X1 p9_mult_21_U552 ( .A1(p9_mult_21_n1021), .A2(p9_mult_21_n1023), 
        .ZN(p9_mult_21_n1045) );
  OAI22_X1 p9_mult_21_U554 ( .A1(p9_mult_21_n911), .A2(p9_mult_21_n1012), .B1(
        p9_mult_21_n903), .B2(p9_mult_21_n1047), .ZN(p9_mult_21_n1018) );
  OAI22_X1 p9_mult_21_U582 ( .A1(p9_mult_21_n905), .A2(p9_mult_21_n1025), .B1(
        B3[6]), .B2(reg4_reg[11]), .ZN(p9_mult_21_n1047) );
  AOI22_X1 p9_mult_21_U555 ( .A1(reg4_reg[11]), .A2(p9_mult_21_n983), .B1(
        B3[7]), .B2(p9_mult_21_n905), .ZN(p9_mult_21_n1012) );
  OAI22_X1 p9_mult_21_U575 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n921), .B1(
        B3[10]), .B2(reg4_reg[7]), .ZN(p9_mult_21_n1042) );
  AOI22_X1 p9_mult_21_U550 ( .A1(B3[11]), .A2(p9_mult_21_n987), .B1(
        reg4_reg[7]), .B2(p9_mult_21_n897), .ZN(p9_mult_21_n1015) );
  OAI21_X1 p9_mult_21_U454 ( .B1(p9_mult_21_n902), .B2(p9_mult_21_n903), .A(
        p9_mult_21_n904), .ZN(p9_mult_21_n874) );
  NAND2_X1 p9_mult_21_U455 ( .A1(p9_mult_21_n880), .A2(p9_mult_21_n882), .ZN(
        p9_mult_21_n904) );
  AOI22_X1 p9_mult_21_U456 ( .A1(B3[13]), .A2(reg4_reg[11]), .B1(
        p9_mult_21_n905), .B2(p9_mult_21_n868), .ZN(p9_mult_21_n882) );
  AOI22_X1 p9_mult_21_U461 ( .A1(reg4_reg[11]), .A2(p9_mult_21_n879), .B1(
        B3[12]), .B2(p9_mult_21_n905), .ZN(p9_mult_21_n902) );
  AOI22_X1 p9_mult_21_U450 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n878), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n896), .ZN(p9_mult_21_n887) );
  OAI22_X1 p9_mult_21_U451 ( .A1(p9_mult_21_n867), .A2(B3[11]), .B1(
        p9_mult_21_n897), .B2(reg4_reg[13]), .ZN(p9_mult_21_n878) );
  AOI222_X1 p9_mult_21_U452 ( .A1(p9_mult_21_n898), .A2(p9_mult_21_n899), .B1(
        p9_mult_21_n898), .B2(p9_mult_21_n900), .C1(p9_mult_21_n899), .C2(
        p9_mult_21_n900), .ZN(p9_mult_21_n886) );
  OAI21_X1 p9_mult_21_U476 ( .B1(p9_mult_21_n936), .B2(p9_mult_21_n937), .A(
        p9_mult_21_n938), .ZN(p9_mult_21_n900) );
  NAND2_X1 p9_mult_21_U477 ( .A1(p9_mult_21_n917), .A2(p9_mult_21_n919), .ZN(
        p9_mult_21_n938) );
  AOI22_X1 p9_mult_21_U497 ( .A1(B3[12]), .A2(p9_mult_21_n939), .B1(
        reg4_reg[9]), .B2(p9_mult_21_n879), .ZN(p9_mult_21_n936) );
  AOI22_X1 p9_mult_21_U466 ( .A1(p9_mult_21_n862), .A2(p9_mult_21_n896), .B1(
        p9_mult_21_n863), .B2(p9_mult_21_n920), .ZN(p9_mult_21_n901) );
  OAI22_X1 p9_mult_21_U475 ( .A1(p9_mult_21_n867), .A2(B3[9]), .B1(
        p9_mult_21_n935), .B2(reg4_reg[13]), .ZN(p9_mult_21_n920) );
  OAI221_X1 p9_mult_21_U830 ( .B1(p9_mult_21_n1379), .B2(p9_mult_21_n867), 
        .C1(reg4_reg[12]), .C2(reg4_reg[13]), .A(p9_mult_21_n1063), .ZN(
        p9_mult_21_n1092) );
  OAI22_X1 p9_mult_21_U467 ( .A1(p9_mult_21_n867), .A2(B3[10]), .B1(
        p9_mult_21_n921), .B2(reg4_reg[13]), .ZN(p9_mult_21_n896) );
  OAI22_X1 p9_mult_21_U888 ( .A1(p9_mult_21_n1379), .A2(p9_mult_21_n905), .B1(
        reg4_reg[11]), .B2(reg4_reg[12]), .ZN(p9_mult_21_n1063) );
  OAI21_X1 p9_mult_21_U464 ( .B1(p9_mult_21_n917), .B2(p9_mult_21_n918), .A(
        p9_mult_21_n919), .ZN(p9_mult_21_n898) );
  AOI22_X1 p9_mult_21_U478 ( .A1(B3[13]), .A2(reg4_reg[9]), .B1(
        p9_mult_21_n939), .B2(p9_mult_21_n868), .ZN(p9_mult_21_n919) );
  XOR2_X1 p9_mult_21_U984 ( .A(p9_mult_21_n1380), .B(p9_mult_21_n1381), .Z(
        p9_mult_21_n1396) );
  XOR2_X1 p9_mult_21_U983 ( .A(p9_mult_21_n1382), .B(p9_mult_21_n1396), .Z(
        p9_mult_21_n1351) );
  XOR2_X1 p9_mult_21_U982 ( .A(p9_mult_21_n1386), .B(p9_mult_21_n1384), .Z(
        p9_mult_21_n1392) );
  XOR2_X1 p9_mult_21_U981 ( .A(p9_mult_21_n1366), .B(p9_mult_21_n1365), .Z(
        p9_mult_21_n1327) );
  XOR2_X1 p9_mult_21_U980 ( .A(p9_mult_21_n1144), .B(p9_mult_21_n1146), .Z(
        p9_mult_21_n1358) );
  XOR2_X1 p9_mult_21_U979 ( .A(p9_mult_21_n1153), .B(p9_mult_21_n1152), .Z(
        p9_mult_21_n1372) );
  XOR2_X1 p9_mult_21_U978 ( .A(p9_mult_21_n1367), .B(p9_mult_21_n1158), .Z(
        p9_mult_21_n1161) );
  XOR2_X1 p9_mult_21_U977 ( .A(p9_mult_21_n1358), .B(p9_mult_21_n1145), .Z(
        p9_mult_21_n1143) );
  XOR2_X1 p9_mult_21_U976 ( .A(p9_mult_21_n1356), .B(p9_mult_21_n1357), .Z(
        p9_mult_21_n1355) );
  XOR2_X1 p9_mult_21_U975 ( .A(p9_mult_21_n1354), .B(p9_mult_21_n1355), .Z(
        p9_mult_21_n1183) );
  XOR2_X1 p9_mult_21_U974 ( .A(p9_mult_21_n1352), .B(p9_mult_21_n1353), .Z(
        p9_mult_21_n1350) );
  XOR2_X1 p9_mult_21_U973 ( .A(p9_mult_21_n1341), .B(p9_mult_21_n1342), .Z(
        p9_mult_21_n1323) );
  XOR2_X1 p9_mult_21_U972 ( .A(p9_mult_21_n1326), .B(p9_mult_21_n1327), .Z(
        p9_mult_21_n1187) );
  XOR2_X1 p9_mult_21_U971 ( .A(p9_mult_21_n1185), .B(p9_mult_21_n1187), .Z(
        p9_mult_21_n1321) );
  XOR2_X1 p9_mult_21_U970 ( .A(p9_mult_21_n1321), .B(p9_mult_21_n1186), .Z(
        p9_mult_21_n1188) );
  XOR2_X1 p9_mult_21_U969 ( .A(p9_mult_21_n1312), .B(p9_mult_21_n1313), .Z(
        p9_mult_21_n1210) );
  XOR2_X1 p9_mult_21_U968 ( .A(p9_mult_21_n1307), .B(p9_mult_21_n1308), .Z(
        p9_mult_21_n1207) );
  XOR2_X1 p9_mult_21_U967 ( .A(p9_mult_21_n1209), .B(p9_mult_21_n1207), .Z(
        p9_mult_21_n1305) );
  XOR2_X1 p9_mult_21_U965 ( .A(p9_mult_21_n1260), .B(p9_mult_21_n1261), .Z(
        p9_mult_21_n1259) );
  XOR2_X1 p9_mult_21_U964 ( .A(p9_mult_21_n1258), .B(p9_mult_21_n1259), .Z(
        p9_mult_21_n1257) );
  XOR2_X1 p9_mult_21_U963 ( .A(p9_mult_21_n1235), .B(p9_mult_21_n1237), .Z(
        p9_mult_21_n1241) );
  XOR2_X1 p9_mult_21_U962 ( .A(p9_mult_21_n1242), .B(p9_mult_21_n1233), .Z(
        p9_mult_21_n1236) );
  XOR2_X1 p9_mult_21_U961 ( .A(p9_mult_21_n1241), .B(p9_mult_21_n1236), .Z(
        p9_mult_21_n1240) );
  XOR2_X1 p9_mult_21_U960 ( .A(p9_mult_21_n1230), .B(p9_mult_21_n1231), .Z(
        p9_mult_21_n1229) );
  XOR2_X1 p9_mult_21_U959 ( .A(p9_mult_21_n1228), .B(p9_mult_21_n1229), .Z(
        p9_mult_21_n1216) );
  XOR2_X1 p9_mult_21_U958 ( .A(p9_mult_21_n1223), .B(p9_mult_21_n1217), .Z(
        p9_mult_21_n1222) );
  XOR2_X1 p9_mult_21_U957 ( .A(p9_mult_21_n1194), .B(p9_mult_21_n1192), .Z(
        p9_mult_21_n1198) );
  XOR2_X1 p9_mult_21_U956 ( .A(p9_mult_21_n1201), .B(p9_mult_21_n1202), .Z(
        p9_mult_21_n1200) );
  XOR2_X1 p9_mult_21_U955 ( .A(p9_mult_21_n1199), .B(p9_mult_21_n1200), .Z(
        p9_mult_21_n1193) );
  XOR2_X1 p9_mult_21_U954 ( .A(n764), .B(p9_mult_21_n1142), .Z(
        p9_mult_21_n1177) );
  XOR2_X1 p9_mult_21_U953 ( .A(p9_mult_21_n1129), .B(p9_mult_21_n1128), .Z(
        p9_mult_21_n1171) );
  XOR2_X1 p9_mult_21_U952 ( .A(p9_mult_21_n1130), .B(p9_mult_21_n1171), .Z(
        p9_mult_21_n1131) );
  XOR2_X1 p9_mult_21_U951 ( .A(p9_mult_21_n1127), .B(p9_mult_21_n1126), .Z(
        p9_mult_21_n1163) );
  XOR2_X1 p9_mult_21_U950 ( .A(p9_mult_21_n1125), .B(p9_mult_21_n1163), .Z(
        p9_mult_21_n1133) );
  XOR2_X1 p9_mult_21_U949 ( .A(p9_mult_21_n1107), .B(p9_mult_21_n1109), .Z(
        p9_mult_21_n1148) );
  XOR2_X1 p9_mult_21_U948 ( .A(p9_mult_21_n1108), .B(p9_mult_21_n1148), .Z(
        p9_mult_21_n1135) );
  XOR2_X1 p9_mult_21_U947 ( .A(p9_mult_21_n1136), .B(p9_mult_21_n1135), .Z(
        p9_mult_21_n1147) );
  XOR2_X1 p9_mult_21_U946 ( .A(p9_mult_21_n1134), .B(p9_mult_21_n1147), .Z(
        p9_mult_21_n1137) );
  XOR2_X1 p9_mult_21_U945 ( .A(p9_mult_21_n1117), .B(p9_mult_21_n1073), .Z(
        p9_mult_21_n1079) );
  XOR2_X1 p9_mult_21_U944 ( .A(p9_mult_21_n1066), .B(p9_mult_21_n1074), .Z(
        p9_mult_21_n1110) );
  XOR2_X1 p9_mult_21_U943 ( .A(p9_mult_21_n1075), .B(p9_mult_21_n1110), .Z(
        p9_mult_21_n1078) );
  XOR2_X1 p9_mult_21_U942 ( .A(p9_mult_21_n1078), .B(p9_mult_21_n1077), .Z(
        p9_mult_21_n1106) );
  XOR2_X1 p9_mult_21_U941 ( .A(p9_mult_21_n1079), .B(p9_mult_21_n1106), .Z(
        p9_mult_21_n1103) );
  XOR2_X1 p9_mult_21_U940 ( .A(p9_mult_21_n1098), .B(p9_mult_21_n1099), .Z(
        p9_mult_21_n1104) );
  XOR2_X1 p9_mult_21_U939 ( .A(p9_mult_21_n1066), .B(p9_mult_21_n1065), .Z(
        p9_mult_21_n1088) );
  XOR2_X1 p9_mult_21_U938 ( .A(p9_mult_21_n1088), .B(p9_mult_21_n1064), .Z(
        p9_mult_21_n1055) );
  XOR2_X1 p9_mult_21_U937 ( .A(p9_mult_21_n1048), .B(p9_mult_21_n1049), .Z(
        p9_mult_21_n1081) );
  XOR2_X1 p9_mult_21_U936 ( .A(p9_mult_21_n1050), .B(p9_mult_21_n1081), .Z(
        p9_mult_21_n1056) );
  XOR2_X1 p9_mult_21_U935 ( .A(p9_mult_21_n1055), .B(p9_mult_21_n1056), .Z(
        p9_mult_21_n1080) );
  XOR2_X1 p9_mult_21_U934 ( .A(p9_mult_21_n1054), .B(p9_mult_21_n1080), .Z(
        p9_mult_21_n1038) );
  XOR2_X1 p9_mult_21_U933 ( .A(p9_mult_21_n1051), .B(p9_mult_21_n1052), .Z(
        p9_mult_21_n1069) );
  XOR2_X1 p9_mult_21_U932 ( .A(p9_mult_21_n1053), .B(p9_mult_21_n1069), .Z(
        p9_mult_21_n1037) );
  XOR2_X1 p9_mult_21_U931 ( .A(p9_mult_21_n1036), .B(p9_mult_21_n1037), .Z(
        p9_mult_21_n1068) );
  XOR2_X1 p9_mult_21_U930 ( .A(p9_mult_21_n1038), .B(p9_mult_21_n1068), .Z(
        p9_mult_21_n1035) );
  XOR2_X1 p9_mult_21_U929 ( .A(p9_mult_21_n1029), .B(p9_mult_21_n1031), .Z(
        p9_mult_21_n1039) );
  XOR2_X1 p9_mult_21_U928 ( .A(p9_mult_21_n1030), .B(p9_mult_21_n1039), .Z(
        p9_mult_21_n1028) );
  XOR2_X1 p9_mult_21_U927 ( .A(p9_mult_21_n1026), .B(p9_mult_21_n1027), .Z(
        p9_mult_21_n1032) );
  XOR2_X1 p9_mult_21_U926 ( .A(p9_mult_21_n1020), .B(p9_mult_21_n991), .Z(
        p9_mult_21_n1001) );
  XOR2_X1 p9_mult_21_U925 ( .A(p9_mult_21_n997), .B(p9_mult_21_n1011), .Z(
        p9_mult_21_n1000) );
  XOR2_X1 p9_mult_21_U924 ( .A(p9_mult_21_n999), .B(p9_mult_21_n1000), .Z(
        p9_mult_21_n1010) );
  XOR2_X1 p9_mult_21_U923 ( .A(p9_mult_21_n1001), .B(p9_mult_21_n1010), .Z(
        p9_mult_21_n979) );
  XOR2_X1 p9_mult_21_U922 ( .A(p9_mult_21_n977), .B(p9_mult_21_n978), .Z(
        p9_mult_21_n1003) );
  XOR2_X1 p9_mult_21_U920 ( .A(p9_mult_21_n946), .B(p9_mult_21_n961), .Z(
        p9_mult_21_n981) );
  XOR2_X1 p9_mult_21_U919 ( .A(p9_mult_21_n967), .B(n774), .Z(p9_mult_21_n973)
         );
  XOR2_X1 p9_mult_21_U918 ( .A(p9_mult_21_n941), .B(p9_mult_21_n942), .Z(
        p9_mult_21_n959) );
  XOR2_X1 p9_mult_21_U917 ( .A(p9_mult_21_n943), .B(p9_mult_21_n959), .Z(
        p9_mult_21_n931) );
  XOR2_X1 p9_mult_21_U916 ( .A(p9_mult_21_n950), .B(p9_mult_21_n944), .Z(
        p9_mult_21_n930) );
  XOR2_X1 p9_mult_21_U915 ( .A(p9_mult_21_n929), .B(p9_mult_21_n930), .Z(
        p9_mult_21_n949) );
  XOR2_X1 p9_mult_21_U914 ( .A(p9_mult_21_n931), .B(p9_mult_21_n949), .Z(
        p9_mult_21_n928) );
  XOR2_X1 p9_mult_21_U913 ( .A(p9_mult_21_n900), .B(p9_mult_21_n913), .Z(
        p9_mult_21_n933) );
  XOR2_X1 p9_mult_21_U912 ( .A(p9_mult_21_n907), .B(p9_mult_21_n908), .Z(
        p9_mult_21_n925) );
  XOR2_X1 p9_mult_21_U911 ( .A(p9_mult_21_n916), .B(p9_mult_21_n898), .Z(
        p9_mult_21_n894) );
  XOR2_X1 p9_mult_21_U910 ( .A(p9_mult_21_n892), .B(p9_mult_21_n893), .Z(
        p9_mult_21_n910) );
  XOR2_X1 p9_mult_21_U909 ( .A(p9_mult_21_n894), .B(p9_mult_21_n910), .Z(
        p9_mult_21_n890) );
  XOR2_X1 p9_mult_21_U908 ( .A(p9_mult_21_n874), .B(p9_mult_21_n886), .Z(
        p9_mult_21_n895) );
  XOR2_X1 p9_mult_21_U906 ( .A(n760), .B(p9_mult_21_n883), .Z(p9_mult_21_n888)
         );
  MUX2_X1 p9_mult_21_U899 ( .A(p9_mult_21_n844), .B(p9_mult_21_n845), .S(
        reg4_reg[0]), .Z(p9_mult_21_n1254) );
  MUX2_X1 p9_mult_21_U897 ( .A(p9_mult_21_n840), .B(p9_mult_21_n841), .S(
        reg4_reg[0]), .Z(p9_mult_21_n1278) );
  MUX2_X1 p9_mult_21_U896 ( .A(p9_mult_21_n838), .B(p9_mult_21_n839), .S(
        reg4_reg[0]), .Z(p9_mult_21_n1270) );
  INV_X1 p11_mult_21_U718 ( .A(p11_mult_21_n267), .ZN(p11_mult_21_n828) );
  INV_X1 p11_mult_21_U719 ( .A(p11_mult_21_n258), .ZN(p11_mult_21_n827) );
  AND3_X1 p11_mult_21_U413 ( .A1(p11_mult_21_n679), .A2(p11_mult_21_n680), 
        .A3(p11_mult_21_n681), .ZN(p11_mult_21_n826) );
  INV_X1 p11_mult_21_U721 ( .A(p11_mult_21_n285), .ZN(p11_mult_21_n832) );
  INV_X1 p11_mult_21_U722 ( .A(p11_mult_21_n278), .ZN(p11_mult_21_n831) );
  AND3_X1 p11_mult_21_U412 ( .A1(p11_mult_21_n660), .A2(p11_mult_21_n661), 
        .A3(p11_mult_21_n662), .ZN(p11_mult_21_n830) );
  OR3_X1 p11_mult_21_U663 ( .A1(p11_mult_21_n741), .A2(A1[0]), .A3(n885), .ZN(
        p11_mult_21_n811) );
  INV_X1 p11_mult_21_U736 ( .A(p11_mult_21_n843), .ZN(p11_mult_21_n845) );
  INV_X1 p11_mult_21_U730 ( .A(A1[0]), .ZN(p11_mult_21_n723) );
  OR2_X1 p11_mult_21_U671 ( .A1(p11_mult_21_n818), .A2(p11_mult_21_n819), .ZN(
        p11_mult_21_n243) );
  INV_X1 p11_mult_21_U503 ( .A(p11_mult_21_n704), .ZN(p11_mult_21_n408) );
  INV_X1 p11_mult_21_U530 ( .A(p11_mult_21_n721), .ZN(p11_mult_21_n394) );
  INV_X1 p11_mult_21_U678 ( .A(p11_mult_21_n231), .ZN(p11_mult_21_n232) );
  INV_X1 p11_mult_21_U423 ( .A(p11_mult_21_n838), .ZN(p11_mult_21_n708) );
  INV_X1 p11_mult_21_U682 ( .A(p11_mult_21_n209), .ZN(p11_mult_21_n210) );
  INV_X1 p11_mult_21_U554 ( .A(p11_mult_21_n739), .ZN(p11_mult_21_n380) );
  INV_X1 p11_mult_21_U687 ( .A(p11_mult_21_n191), .ZN(p11_mult_21_n192) );
  INV_X1 p11_mult_21_U581 ( .A(p11_mult_21_n756), .ZN(p11_mult_21_n366) );
  NAND2_X1 p11_mult_21_U690 ( .A1(p11_mult_21_n741), .A2(p11_mult_21_n822), 
        .ZN(p11_mult_21_n743) );
  INV_X1 p11_mult_21_U694 ( .A(p11_mult_21_n177), .ZN(p11_mult_21_n178) );
  INV_X1 p11_mult_21_U608 ( .A(p11_mult_21_n773), .ZN(p11_mult_21_n352) );
  INV_X1 p11_mult_21_U701 ( .A(p11_mult_21_n167), .ZN(p11_mult_21_n168) );
  INV_X1 p11_mult_21_U710 ( .A(p11_mult_21_n792), .ZN(p11_mult_21_n688) );
  INV_X1 p11_mult_21_U711 ( .A(p11_mult_21_n794), .ZN(p11_mult_21_n687) );
  INV_X1 p11_mult_21_U632 ( .A(p11_mult_21_n790), .ZN(p11_mult_21_n338) );
  INV_X1 p11_mult_21_U658 ( .A(p11_mult_21_n807), .ZN(p11_mult_21_n806) );
  NAND2_X1 p11_mult_21_U697 ( .A1(p11_mult_21_n758), .A2(p11_mult_21_n823), 
        .ZN(p11_mult_21_n760) );
  NAND2_X1 p11_mult_21_U704 ( .A1(p11_mult_21_n775), .A2(p11_mult_21_n824), 
        .ZN(p11_mult_21_n777) );
  NAND2_X1 p11_mult_21_U725 ( .A1(p11_mult_21_n708), .A2(p11_mult_21_n839), 
        .ZN(p11_mult_21_n707) );
  NAND2_X1 p11_mult_21_U475 ( .A1(p11_mult_21_n724), .A2(p11_mult_21_n820), 
        .ZN(p11_mult_21_n726) );
  NAND2_X1 p11_mult_21_U712 ( .A1(p11_mult_21_n792), .A2(p11_mult_21_n825), 
        .ZN(p11_mult_21_n794) );
  NAND2_X1 p11_mult_21_U459 ( .A1(p11_mult_21_n234), .A2(p11_mult_21_n245), 
        .ZN(p11_mult_21_n671) );
  NAND2_X1 p11_mult_21_U472 ( .A1(p11_mult_21_n277), .A2(p11_mult_21_n268), 
        .ZN(p11_mult_21_n681) );
  OAI22_X1 p11_mult_21_U565 ( .A1(p11_mult_21_n747), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n748), .ZN(p11_mult_21_n374) );
  OAI222_X1 p11_mult_21_U720 ( .A1(p11_mult_21_n830), .A2(p11_mult_21_n831), 
        .B1(p11_mult_21_n830), .B2(p11_mult_21_n832), .C1(p11_mult_21_n832), 
        .C2(p11_mult_21_n831), .ZN(p11_mult_21_n829) );
  OAI22_X1 p11_mult_21_U495 ( .A1(p11_mult_21_n699), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n700), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n412) );
  NOR2_X1 p11_mult_21_U610 ( .A1(p11_mult_21_n723), .A2(p11_mult_21_n775), 
        .ZN(p11_mult_21_n351) );
  OAI22_X1 p11_mult_21_U563 ( .A1(p11_mult_21_n746), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n747), .ZN(p11_mult_21_n375) );
  XNOR2_X1 p11_mult_21_U566 ( .A(A1[4]), .B(reg2[7]), .ZN(p11_mult_21_n747) );
  OAI22_X1 p11_mult_21_U543 ( .A1(p11_mult_21_n731), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n732), .ZN(p11_mult_21_n387) );
  XNOR2_X1 p11_mult_21_U523 ( .A(A1[8]), .B(reg2[3]), .ZN(p11_mult_21_n716) );
  OAI22_X1 p11_mult_21_U586 ( .A1(p11_mult_21_n761), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n762), .ZN(p11_mult_21_n363) );
  NAND2_X1 p11_mult_21_U447 ( .A1(p11_mult_21_n293), .A2(p11_mult_21_n286), 
        .ZN(p11_mult_21_n662) );
  NAND2_X1 p11_mult_21_U446 ( .A1(p11_mult_21_n635), .A2(p11_mult_21_n293), 
        .ZN(p11_mult_21_n661) );
  NAND2_X1 p11_mult_21_U445 ( .A1(p11_mult_21_n635), .A2(p11_mult_21_n286), 
        .ZN(p11_mult_21_n660) );
  OAI22_X1 p11_mult_21_U493 ( .A1(p11_mult_21_n698), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n699), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n413) );
  XNOR2_X1 p11_mult_21_U587 ( .A(A1[1]), .B(reg2[9]), .ZN(p11_mult_21_n761) );
  XNOR2_X1 p11_mult_21_U521 ( .A(A1[7]), .B(reg2[3]), .ZN(p11_mult_21_n715) );
  OAI22_X1 p11_mult_21_U541 ( .A1(p11_mult_21_n730), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n731), .ZN(p11_mult_21_n388) );
  XNOR2_X1 p11_mult_21_U544 ( .A(A1[5]), .B(reg2[5]), .ZN(p11_mult_21_n731) );
  OAI22_X1 p11_mult_21_U561 ( .A1(p11_mult_21_n745), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n746), .ZN(p11_mult_21_n376) );
  XNOR2_X1 p11_mult_21_U564 ( .A(A1[3]), .B(reg2[7]), .ZN(p11_mult_21_n746) );
  NAND2_X1 p11_mult_21_U418 ( .A1(p11_mult_21_n299), .A2(p11_mult_21_n294), 
        .ZN(p11_mult_21_n642) );
  XNOR2_X1 p11_mult_21_U519 ( .A(A1[6]), .B(reg2[3]), .ZN(p11_mult_21_n714) );
  OAI22_X1 p11_mult_21_U559 ( .A1(p11_mult_21_n744), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n745), .ZN(p11_mult_21_n377) );
  XNOR2_X1 p11_mult_21_U562 ( .A(A1[2]), .B(reg2[7]), .ZN(p11_mult_21_n745) );
  OAI22_X1 p11_mult_21_U491 ( .A1(p11_mult_21_n697), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n698), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n414) );
  NOR2_X1 p11_mult_21_U583 ( .A1(p11_mult_21_n723), .A2(p11_mult_21_n758), 
        .ZN(p11_mult_21_n365) );
  OAI22_X1 p11_mult_21_U539 ( .A1(p11_mult_21_n729), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n730), .ZN(p11_mult_21_n389) );
  XNOR2_X1 p11_mult_21_U542 ( .A(A1[4]), .B(reg2[5]), .ZN(p11_mult_21_n730) );
  XNOR2_X1 p11_mult_21_U517 ( .A(A1[5]), .B(reg2[3]), .ZN(p11_mult_21_n713) );
  OAI22_X1 p11_mult_21_U489 ( .A1(p11_mult_21_n696), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n697), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n415) );
  OAI22_X1 p11_mult_21_U537 ( .A1(p11_mult_21_n728), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n729), .ZN(p11_mult_21_n390) );
  XNOR2_X1 p11_mult_21_U540 ( .A(A1[3]), .B(reg2[5]), .ZN(p11_mult_21_n729) );
  OAI22_X1 p11_mult_21_U557 ( .A1(p11_mult_21_n742), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n744), .ZN(p11_mult_21_n378) );
  XNOR2_X1 p11_mult_21_U560 ( .A(A1[1]), .B(reg2[7]), .ZN(p11_mult_21_n744) );
  XNOR2_X1 p11_mult_21_U558 ( .A(reg2[7]), .B(A1[0]), .ZN(p11_mult_21_n742) );
  OAI21_X1 p11_mult_21_U662 ( .B1(n885), .B2(p11_mult_21_n743), .A(
        p11_mult_21_n811), .ZN(p11_mult_21_n320) );
  XNOR2_X1 p11_mult_21_U515 ( .A(A1[4]), .B(reg2[3]), .ZN(p11_mult_21_n712) );
  NOR2_X1 p11_mult_21_U556 ( .A1(p11_mult_21_n723), .A2(p11_mult_21_n741), 
        .ZN(p11_mult_21_n379) );
  OAI22_X1 p11_mult_21_U487 ( .A1(p11_mult_21_n695), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n696), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n416) );
  XNOR2_X1 p11_mult_21_U538 ( .A(A1[2]), .B(reg2[5]), .ZN(p11_mult_21_n728) );
  XNOR2_X1 p11_mult_21_U536 ( .A(A1[1]), .B(reg2[5]), .ZN(p11_mult_21_n727) );
  OAI22_X1 p11_mult_21_U485 ( .A1(p11_mult_21_n694), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n695), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n417) );
  XNOR2_X1 p11_mult_21_U513 ( .A(A1[3]), .B(reg2[3]), .ZN(p11_mult_21_n711) );
  XNOR2_X1 p11_mult_21_U511 ( .A(A1[2]), .B(reg2[3]), .ZN(p11_mult_21_n710) );
  NOR2_X1 p11_mult_21_U532 ( .A1(p11_mult_21_n723), .A2(p11_mult_21_n724), 
        .ZN(p11_mult_21_n393) );
  OAI22_X1 p11_mult_21_U483 ( .A1(p11_mult_21_n692), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n694), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n418) );
  XNOR2_X1 p11_mult_21_U509 ( .A(A1[1]), .B(reg2[3]), .ZN(p11_mult_21_n709) );
  XNOR2_X1 p11_mult_21_U507 ( .A(reg2[3]), .B(A1[0]), .ZN(p11_mult_21_n706) );
  NAND2_X1 p11_mult_21_U731 ( .A1(p11_mult_21_n843), .A2(p11_mult_21_n844), 
        .ZN(p11_mult_21_n842) );
  NAND2_X1 p11_mult_21_U732 ( .A1(p11_mult_21_n844), .A2(p11_mult_21_n838), 
        .ZN(p11_mult_21_n841) );
  OAI22_X1 p11_mult_21_U733 ( .A1(p11_mult_21_n845), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n690), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n844) );
  NOR2_X1 p11_mult_21_U737 ( .A1(n888), .A2(A1[1]), .ZN(p11_mult_21_n843) );
  OAI22_X1 p11_mult_21_U497 ( .A1(p11_mult_21_n700), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n701), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n411) );
  OAI22_X1 p11_mult_21_U545 ( .A1(p11_mult_21_n732), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n733), .ZN(p11_mult_21_n386) );
  XNOR2_X1 p11_mult_21_U546 ( .A(A1[6]), .B(reg2[5]), .ZN(p11_mult_21_n732) );
  OAI22_X1 p11_mult_21_U588 ( .A1(p11_mult_21_n762), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n763), .ZN(p11_mult_21_n362) );
  XNOR2_X1 p11_mult_21_U589 ( .A(A1[2]), .B(reg2[9]), .ZN(p11_mult_21_n762) );
  OAI22_X1 p11_mult_21_U547 ( .A1(p11_mult_21_n733), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n734), .ZN(p11_mult_21_n385) );
  XNOR2_X1 p11_mult_21_U548 ( .A(A1[7]), .B(reg2[5]), .ZN(p11_mult_21_n733) );
  OAI22_X1 p11_mult_21_U567 ( .A1(p11_mult_21_n748), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n749), .ZN(p11_mult_21_n373) );
  XNOR2_X1 p11_mult_21_U568 ( .A(A1[5]), .B(reg2[7]), .ZN(p11_mult_21_n748) );
  XNOR2_X1 p11_mult_21_U525 ( .A(A1[9]), .B(reg2[3]), .ZN(p11_mult_21_n717) );
  OAI22_X1 p11_mult_21_U613 ( .A1(p11_mult_21_n778), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n779), .ZN(p11_mult_21_n349) );
  XNOR2_X1 p11_mult_21_U614 ( .A(A1[1]), .B(reg2[11]), .ZN(p11_mult_21_n778)
         );
  OAI22_X1 p11_mult_21_U499 ( .A1(p11_mult_21_n701), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n702), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n410) );
  NOR2_X1 p11_mult_21_U634 ( .A1(p11_mult_21_n723), .A2(p11_mult_21_n792), 
        .ZN(p11_mult_21_n337) );
  OAI22_X1 p11_mult_21_U590 ( .A1(p11_mult_21_n763), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n764), .ZN(p11_mult_21_n361) );
  XNOR2_X1 p11_mult_21_U591 ( .A(A1[3]), .B(reg2[9]), .ZN(p11_mult_21_n763) );
  OAI22_X1 p11_mult_21_U592 ( .A1(p11_mult_21_n764), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n765), .ZN(p11_mult_21_n360) );
  XNOR2_X1 p11_mult_21_U593 ( .A(A1[4]), .B(reg2[9]), .ZN(p11_mult_21_n764) );
  OAI22_X1 p11_mult_21_U549 ( .A1(p11_mult_21_n734), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n735), .ZN(p11_mult_21_n384) );
  XNOR2_X1 p11_mult_21_U550 ( .A(A1[8]), .B(reg2[5]), .ZN(p11_mult_21_n734) );
  OAI22_X1 p11_mult_21_U615 ( .A1(p11_mult_21_n779), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n780), .ZN(p11_mult_21_n348) );
  XNOR2_X1 p11_mult_21_U616 ( .A(A1[2]), .B(reg2[11]), .ZN(p11_mult_21_n779)
         );
  XNOR2_X1 p11_mult_21_U670 ( .A(p11_mult_21_n818), .B(p11_mult_21_n819), .ZN(
        p11_mult_21_n244) );
  XNOR2_X1 p11_mult_21_U527 ( .A(A1[10]), .B(reg2[3]), .ZN(p11_mult_21_n718)
         );
  OAI22_X1 p11_mult_21_U569 ( .A1(p11_mult_21_n749), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n750), .ZN(p11_mult_21_n372) );
  XNOR2_X1 p11_mult_21_U570 ( .A(A1[6]), .B(reg2[7]), .ZN(p11_mult_21_n749) );
  OAI22_X1 p11_mult_21_U501 ( .A1(p11_mult_21_n702), .A2(p11_mult_21_n691), 
        .B1(p11_mult_21_n703), .B2(p11_mult_21_n693), .ZN(p11_mult_21_n409) );
  OAI22_X1 p11_mult_21_U635 ( .A1(p11_mult_21_n793), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n795), .ZN(p11_mult_21_n336) );
  XNOR2_X1 p11_mult_21_U636 ( .A(reg2[13]), .B(A1[0]), .ZN(p11_mult_21_n793)
         );
  OAI21_X1 p11_mult_21_U668 ( .B1(n887), .B2(p11_mult_21_n794), .A(
        p11_mult_21_n817), .ZN(p11_mult_21_n317) );
  OAI22_X1 p11_mult_21_U571 ( .A1(p11_mult_21_n750), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n751), .ZN(p11_mult_21_n371) );
  XNOR2_X1 p11_mult_21_U572 ( .A(A1[7]), .B(reg2[7]), .ZN(p11_mult_21_n750) );
  OAI22_X1 p11_mult_21_U637 ( .A1(p11_mult_21_n795), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n796), .ZN(p11_mult_21_n335) );
  XNOR2_X1 p11_mult_21_U638 ( .A(A1[1]), .B(reg2[13]), .ZN(p11_mult_21_n795)
         );
  OAI22_X1 p11_mult_21_U672 ( .A1(p11_mult_21_n735), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n736), .ZN(p11_mult_21_n819) );
  XNOR2_X1 p11_mult_21_U674 ( .A(A1[9]), .B(reg2[5]), .ZN(p11_mult_21_n735) );
  OAI22_X1 p11_mult_21_U675 ( .A1(p11_mult_21_n780), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n781), .ZN(p11_mult_21_n818) );
  XNOR2_X1 p11_mult_21_U677 ( .A(A1[3]), .B(reg2[11]), .ZN(p11_mult_21_n780)
         );
  AOI21_X1 p11_mult_21_U504 ( .B1(p11_mult_21_n691), .B2(p11_mult_21_n693), 
        .A(p11_mult_21_n703), .ZN(p11_mult_21_n704) );
  OAI22_X1 p11_mult_21_U594 ( .A1(p11_mult_21_n765), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n766), .ZN(p11_mult_21_n359) );
  XNOR2_X1 p11_mult_21_U595 ( .A(A1[5]), .B(reg2[9]), .ZN(p11_mult_21_n765) );
  XNOR2_X1 p11_mult_21_U529 ( .A(A1[11]), .B(reg2[3]), .ZN(p11_mult_21_n719)
         );
  OAI22_X1 p11_mult_21_U641 ( .A1(p11_mult_21_n797), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n798), .ZN(p11_mult_21_n333) );
  OAI22_X1 p11_mult_21_U600 ( .A1(p11_mult_21_n768), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n769), .ZN(p11_mult_21_n356) );
  OAI22_X1 p11_mult_21_U643 ( .A1(p11_mult_21_n798), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n799), .ZN(p11_mult_21_n332) );
  XNOR2_X1 p11_mult_21_U644 ( .A(A1[4]), .B(reg2[13]), .ZN(p11_mult_21_n798)
         );
  OAI22_X1 p11_mult_21_U596 ( .A1(p11_mult_21_n766), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n767), .ZN(p11_mult_21_n358) );
  XNOR2_X1 p11_mult_21_U597 ( .A(A1[6]), .B(reg2[9]), .ZN(p11_mult_21_n766) );
  OAI22_X1 p11_mult_21_U573 ( .A1(p11_mult_21_n751), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n752), .ZN(p11_mult_21_n370) );
  XNOR2_X1 p11_mult_21_U574 ( .A(A1[8]), .B(reg2[7]), .ZN(p11_mult_21_n751) );
  OAI22_X1 p11_mult_21_U639 ( .A1(p11_mult_21_n796), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n797), .ZN(p11_mult_21_n334) );
  XNOR2_X1 p11_mult_21_U642 ( .A(A1[3]), .B(reg2[13]), .ZN(p11_mult_21_n797)
         );
  XNOR2_X1 p11_mult_21_U640 ( .A(A1[2]), .B(reg2[13]), .ZN(p11_mult_21_n796)
         );
  OAI22_X1 p11_mult_21_U575 ( .A1(p11_mult_21_n752), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n753), .ZN(p11_mult_21_n369) );
  XNOR2_X1 p11_mult_21_U576 ( .A(A1[9]), .B(reg2[7]), .ZN(p11_mult_21_n752) );
  XNOR2_X1 p11_mult_21_U680 ( .A(A1[13]), .B(reg2[3]), .ZN(p11_mult_21_n722)
         );
  XNOR2_X1 p11_mult_21_U726 ( .A(n575), .B(reg2[2]), .ZN(p11_mult_21_n839) );
  XNOR2_X1 p11_mult_21_U681 ( .A(A1[12]), .B(reg2[3]), .ZN(p11_mult_21_n720)
         );
  OAI22_X1 p11_mult_21_U617 ( .A1(p11_mult_21_n781), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n782), .ZN(p11_mult_21_n346) );
  XNOR2_X1 p11_mult_21_U676 ( .A(A1[4]), .B(reg2[11]), .ZN(p11_mult_21_n781)
         );
  OAI22_X1 p11_mult_21_U551 ( .A1(p11_mult_21_n736), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n737), .ZN(p11_mult_21_n382) );
  XNOR2_X1 p11_mult_21_U673 ( .A(A1[10]), .B(reg2[5]), .ZN(p11_mult_21_n736)
         );
  OAI22_X1 p11_mult_21_U598 ( .A1(p11_mult_21_n767), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n768), .ZN(p11_mult_21_n357) );
  XNOR2_X1 p11_mult_21_U601 ( .A(A1[8]), .B(reg2[9]), .ZN(p11_mult_21_n768) );
  XNOR2_X1 p11_mult_21_U599 ( .A(A1[7]), .B(reg2[9]), .ZN(p11_mult_21_n767) );
  OAI22_X1 p11_mult_21_U552 ( .A1(p11_mult_21_n737), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n738), .ZN(p11_mult_21_n381) );
  XNOR2_X1 p11_mult_21_U553 ( .A(A1[11]), .B(reg2[5]), .ZN(p11_mult_21_n737)
         );
  OAI22_X1 p11_mult_21_U618 ( .A1(p11_mult_21_n782), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n783), .ZN(p11_mult_21_n345) );
  XNOR2_X1 p11_mult_21_U619 ( .A(A1[5]), .B(reg2[11]), .ZN(p11_mult_21_n782)
         );
  OAI22_X1 p11_mult_21_U620 ( .A1(p11_mult_21_n783), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n784), .ZN(p11_mult_21_n344) );
  XNOR2_X1 p11_mult_21_U621 ( .A(A1[6]), .B(reg2[11]), .ZN(p11_mult_21_n783)
         );
  OAI22_X1 p11_mult_21_U577 ( .A1(p11_mult_21_n753), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n754), .ZN(p11_mult_21_n368) );
  XNOR2_X1 p11_mult_21_U578 ( .A(A1[10]), .B(reg2[7]), .ZN(p11_mult_21_n753)
         );
  OAI22_X1 p11_mult_21_U579 ( .A1(p11_mult_21_n754), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n755), .ZN(p11_mult_21_n367) );
  XNOR2_X1 p11_mult_21_U580 ( .A(A1[11]), .B(reg2[7]), .ZN(p11_mult_21_n754)
         );
  OAI22_X1 p11_mult_21_U622 ( .A1(p11_mult_21_n784), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n785), .ZN(p11_mult_21_n343) );
  XNOR2_X1 p11_mult_21_U623 ( .A(A1[7]), .B(reg2[11]), .ZN(p11_mult_21_n784)
         );
  OAI22_X1 p11_mult_21_U602 ( .A1(p11_mult_21_n769), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n770), .ZN(p11_mult_21_n355) );
  XNOR2_X1 p11_mult_21_U603 ( .A(A1[9]), .B(reg2[9]), .ZN(p11_mult_21_n769) );
  OAI22_X1 p11_mult_21_U604 ( .A1(p11_mult_21_n770), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n771), .ZN(p11_mult_21_n354) );
  XNOR2_X1 p11_mult_21_U605 ( .A(A1[10]), .B(reg2[9]), .ZN(p11_mult_21_n770)
         );
  AOI21_X1 p11_mult_21_U555 ( .B1(p11_mult_21_n726), .B2(p11_mult_21_n724), 
        .A(p11_mult_21_n740), .ZN(p11_mult_21_n739) );
  OAI22_X1 p11_mult_21_U645 ( .A1(p11_mult_21_n799), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n800), .ZN(p11_mult_21_n331) );
  XNOR2_X1 p11_mult_21_U646 ( .A(A1[5]), .B(reg2[13]), .ZN(p11_mult_21_n799)
         );
  OAI22_X1 p11_mult_21_U683 ( .A1(p11_mult_21_n738), .A2(p11_mult_21_n726), 
        .B1(p11_mult_21_n724), .B2(p11_mult_21_n740), .ZN(p11_mult_21_n209) );
  XNOR2_X1 p11_mult_21_U684 ( .A(A1[13]), .B(reg2[5]), .ZN(p11_mult_21_n740)
         );
  XNOR2_X1 p11_mult_21_U685 ( .A(n886), .B(reg2[4]), .ZN(p11_mult_21_n820) );
  XNOR2_X1 p11_mult_21_U686 ( .A(A1[12]), .B(reg2[5]), .ZN(p11_mult_21_n738)
         );
  OAI22_X1 p11_mult_21_U624 ( .A1(p11_mult_21_n785), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n786), .ZN(p11_mult_21_n342) );
  XNOR2_X1 p11_mult_21_U625 ( .A(A1[8]), .B(reg2[11]), .ZN(p11_mult_21_n785)
         );
  OAI22_X1 p11_mult_21_U647 ( .A1(p11_mult_21_n800), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n801), .ZN(p11_mult_21_n330) );
  XNOR2_X1 p11_mult_21_U648 ( .A(A1[6]), .B(reg2[13]), .ZN(p11_mult_21_n800)
         );
  OAI22_X1 p11_mult_21_U606 ( .A1(p11_mult_21_n771), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n772), .ZN(p11_mult_21_n353) );
  XNOR2_X1 p11_mult_21_U607 ( .A(A1[11]), .B(reg2[9]), .ZN(p11_mult_21_n771)
         );
  OAI22_X1 p11_mult_21_U626 ( .A1(p11_mult_21_n786), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n787), .ZN(p11_mult_21_n341) );
  XNOR2_X1 p11_mult_21_U627 ( .A(A1[9]), .B(reg2[11]), .ZN(p11_mult_21_n786)
         );
  AOI21_X1 p11_mult_21_U582 ( .B1(p11_mult_21_n743), .B2(p11_mult_21_n741), 
        .A(p11_mult_21_n757), .ZN(p11_mult_21_n756) );
  OAI22_X1 p11_mult_21_U649 ( .A1(p11_mult_21_n801), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n802), .ZN(p11_mult_21_n329) );
  XNOR2_X1 p11_mult_21_U650 ( .A(A1[7]), .B(reg2[13]), .ZN(p11_mult_21_n801)
         );
  OAI22_X1 p11_mult_21_U688 ( .A1(p11_mult_21_n755), .A2(p11_mult_21_n743), 
        .B1(p11_mult_21_n741), .B2(p11_mult_21_n757), .ZN(p11_mult_21_n191) );
  XNOR2_X1 p11_mult_21_U689 ( .A(A1[13]), .B(reg2[7]), .ZN(p11_mult_21_n757)
         );
  XNOR2_X1 p11_mult_21_U691 ( .A(n885), .B(reg2[6]), .ZN(p11_mult_21_n822) );
  XNOR2_X1 p11_mult_21_U693 ( .A(A1[12]), .B(reg2[7]), .ZN(p11_mult_21_n755)
         );
  OAI22_X1 p11_mult_21_U630 ( .A1(p11_mult_21_n788), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n789), .ZN(p11_mult_21_n339) );
  OAI22_X1 p11_mult_21_U628 ( .A1(p11_mult_21_n787), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n788), .ZN(p11_mult_21_n340) );
  XNOR2_X1 p11_mult_21_U631 ( .A(A1[11]), .B(reg2[11]), .ZN(p11_mult_21_n788)
         );
  XNOR2_X1 p11_mult_21_U629 ( .A(A1[10]), .B(reg2[11]), .ZN(p11_mult_21_n787)
         );
  OAI22_X1 p11_mult_21_U651 ( .A1(p11_mult_21_n802), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n803), .ZN(p11_mult_21_n328) );
  XNOR2_X1 p11_mult_21_U652 ( .A(A1[8]), .B(reg2[13]), .ZN(p11_mult_21_n802)
         );
  AOI21_X1 p11_mult_21_U609 ( .B1(p11_mult_21_n760), .B2(p11_mult_21_n758), 
        .A(p11_mult_21_n774), .ZN(p11_mult_21_n773) );
  OAI22_X1 p11_mult_21_U695 ( .A1(p11_mult_21_n772), .A2(p11_mult_21_n760), 
        .B1(p11_mult_21_n758), .B2(p11_mult_21_n774), .ZN(p11_mult_21_n177) );
  XNOR2_X1 p11_mult_21_U696 ( .A(A1[13]), .B(reg2[9]), .ZN(p11_mult_21_n774)
         );
  XNOR2_X1 p11_mult_21_U698 ( .A(n884), .B(reg2[8]), .ZN(p11_mult_21_n823) );
  XNOR2_X1 p11_mult_21_U700 ( .A(A1[12]), .B(reg2[9]), .ZN(p11_mult_21_n772)
         );
  OAI22_X1 p11_mult_21_U653 ( .A1(p11_mult_21_n803), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n804), .ZN(p11_mult_21_n327) );
  XNOR2_X1 p11_mult_21_U654 ( .A(A1[9]), .B(reg2[13]), .ZN(p11_mult_21_n803)
         );
  OAI22_X1 p11_mult_21_U655 ( .A1(p11_mult_21_n804), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n805), .ZN(p11_mult_21_n326) );
  XNOR2_X1 p11_mult_21_U656 ( .A(A1[10]), .B(reg2[13]), .ZN(p11_mult_21_n804)
         );
  AOI22_X1 p11_mult_21_U708 ( .A1(p11_mult_21_n807), .A2(p11_mult_21_n687), 
        .B1(p11_mult_21_n688), .B2(p11_mult_21_n689), .ZN(p11_mult_21_n162) );
  XNOR2_X1 p11_mult_21_U709 ( .A(A1[13]), .B(n887), .ZN(p11_mult_21_n689) );
  AOI21_X1 p11_mult_21_U633 ( .B1(p11_mult_21_n777), .B2(p11_mult_21_n775), 
        .A(p11_mult_21_n791), .ZN(p11_mult_21_n790) );
  OAI22_X1 p11_mult_21_U702 ( .A1(p11_mult_21_n789), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n775), .B2(p11_mult_21_n791), .ZN(p11_mult_21_n167) );
  XNOR2_X1 p11_mult_21_U703 ( .A(A1[13]), .B(reg2[11]), .ZN(p11_mult_21_n791)
         );
  XNOR2_X1 p11_mult_21_U705 ( .A(n883), .B(reg2[10]), .ZN(p11_mult_21_n824) );
  XNOR2_X1 p11_mult_21_U707 ( .A(A1[12]), .B(reg2[11]), .ZN(p11_mult_21_n789)
         );
  OAI22_X1 p11_mult_21_U657 ( .A1(p11_mult_21_n805), .A2(p11_mult_21_n794), 
        .B1(p11_mult_21_n792), .B2(p11_mult_21_n806), .ZN(p11_mult_21_n325) );
  XNOR2_X1 p11_mult_21_U713 ( .A(n887), .B(reg2[12]), .ZN(p11_mult_21_n825) );
  XNOR2_X1 p11_mult_21_U659 ( .A(A1[11]), .B(reg2[13]), .ZN(p11_mult_21_n805)
         );
  XOR2_X1 p11_mult_21_U739 ( .A(reg2[2]), .B(reg2[1]), .Z(p11_mult_21_n838) );
  MUX2_X1 p11_mult_21_U729 ( .A(p11_mult_21_n841), .B(p11_mult_21_n842), .S(
        p11_mult_21_n723), .Z(p11_mult_21_n840) );
  XOR2_X1 p11_mult_21_U716 ( .A(A1[12]), .B(reg2[13]), .Z(p11_mult_21_n807) );
  NAND3_X1 p11_mult_21_U669 ( .A1(p11_mult_21_n688), .A2(p11_mult_21_n723), 
        .A3(reg2[13]), .ZN(p11_mult_21_n817) );
  XOR2_X1 p11_mult_21_U505 ( .A(A1[13]), .B(n888), .Z(p11_mult_21_n703) );
  XOR2_X1 p11_mult_21_U462 ( .A(p11_mult_21_n659), .B(p11_mult_21_n672), .Z(
        temp6[0]) );
  XOR2_X1 p11_mult_21_U461 ( .A(p11_mult_21_n246), .B(p11_mult_21_n257), .Z(
        p11_mult_21_n672) );
  XOR2_X1 p11_mult_21_U456 ( .A(p11_mult_21_n148), .B(p11_mult_21_n668), .Z(
        temp6[1]) );
  XOR2_X1 p11_mult_21_U455 ( .A(p11_mult_21_n234), .B(p11_mult_21_n245), .Z(
        p11_mult_21_n668) );
  XOR2_X1 p11_mult_21_U436 ( .A(p11_mult_21_n651), .B(p11_mult_21_n652), .Z(
        temp6[2]) );
  XOR2_X1 p11_mult_21_U435 ( .A(p11_mult_21_n222), .B(p11_mult_21_n233), .Z(
        p11_mult_21_n652) );
  NAND3_X1 p11_mult_21_U433 ( .A1(p11_mult_21_n669), .A2(p11_mult_21_n670), 
        .A3(p11_mult_21_n671), .ZN(p11_mult_21_n651) );
  XOR2_X1 p11_mult_21_U428 ( .A(p11_mult_21_n143), .B(p11_mult_21_n646), .Z(
        temp6[6]) );
  XOR2_X1 p11_mult_21_U427 ( .A(p11_mult_21_n193), .B(p11_mult_21_n186), .Z(
        p11_mult_21_n646) );
  NAND3_X1 p11_mult_21_U409 ( .A1(p11_mult_21_n640), .A2(p11_mult_21_n641), 
        .A3(p11_mult_21_n642), .ZN(p11_mult_21_n635) );
  FA_X1 p11_mult_21_U144 ( .A(p11_mult_21_n418), .B(p11_mult_21_n393), .CI(
        p11_mult_21_n405), .CO(p11_mult_21_n313), .S(p11_mult_21_n314) );
  FA_X1 p11_mult_21_U141 ( .A(p11_mult_21_n416), .B(p11_mult_21_n379), .CI(
        p11_mult_21_n403), .CO(p11_mult_21_n307), .S(p11_mult_21_n308) );
  HA_X1 p11_mult_21_U139 ( .A(p11_mult_21_n320), .B(p11_mult_21_n378), .CO(
        p11_mult_21_n303), .S(p11_mult_21_n304) );
  FA_X1 p11_mult_21_U138 ( .A(p11_mult_21_n390), .B(p11_mult_21_n415), .CI(
        p11_mult_21_n402), .CO(p11_mult_21_n301), .S(p11_mult_21_n302) );
  FA_X1 p11_mult_21_U137 ( .A(p11_mult_21_n307), .B(p11_mult_21_n304), .CI(
        p11_mult_21_n302), .CO(p11_mult_21_n299), .S(p11_mult_21_n300) );
  FA_X1 p11_mult_21_U136 ( .A(p11_mult_21_n389), .B(p11_mult_21_n365), .CI(
        p11_mult_21_n414), .CO(p11_mult_21_n297), .S(p11_mult_21_n298) );
  FA_X1 p11_mult_21_U135 ( .A(p11_mult_21_n377), .B(p11_mult_21_n401), .CI(
        p11_mult_21_n303), .CO(p11_mult_21_n295), .S(p11_mult_21_n296) );
  FA_X1 p11_mult_21_U134 ( .A(p11_mult_21_n298), .B(p11_mult_21_n301), .CI(
        p11_mult_21_n296), .CO(p11_mult_21_n293), .S(p11_mult_21_n294) );
  FA_X1 p11_mult_21_U132 ( .A(p11_mult_21_n376), .B(p11_mult_21_n388), .CI(
        p11_mult_21_n400), .CO(p11_mult_21_n289), .S(p11_mult_21_n290) );
  FA_X1 p11_mult_21_U131 ( .A(p11_mult_21_n292), .B(p11_mult_21_n413), .CI(
        p11_mult_21_n297), .CO(p11_mult_21_n287), .S(p11_mult_21_n288) );
  FA_X1 p11_mult_21_U130 ( .A(p11_mult_21_n290), .B(p11_mult_21_n295), .CI(
        p11_mult_21_n288), .CO(p11_mult_21_n285), .S(p11_mult_21_n286) );
  FA_X1 p11_mult_21_U129 ( .A(p11_mult_21_n375), .B(p11_mult_21_n351), .CI(
        p11_mult_21_n412), .CO(p11_mult_21_n283), .S(p11_mult_21_n284) );
  FA_X1 p11_mult_21_U128 ( .A(p11_mult_21_n363), .B(p11_mult_21_n399), .CI(
        p11_mult_21_n387), .CO(p11_mult_21_n281), .S(p11_mult_21_n282) );
  FA_X1 p11_mult_21_U127 ( .A(p11_mult_21_n289), .B(p11_mult_21_n291), .CI(
        p11_mult_21_n284), .CO(p11_mult_21_n279), .S(p11_mult_21_n280) );
  FA_X1 p11_mult_21_U126 ( .A(p11_mult_21_n287), .B(p11_mult_21_n282), .CI(
        p11_mult_21_n280), .CO(p11_mult_21_n277), .S(p11_mult_21_n278) );
  FA_X1 p11_mult_21_U124 ( .A(p11_mult_21_n362), .B(p11_mult_21_n386), .CI(
        p11_mult_21_n411), .CO(p11_mult_21_n273), .S(p11_mult_21_n274) );
  FA_X1 p11_mult_21_U123 ( .A(p11_mult_21_n374), .B(p11_mult_21_n398), .CI(
        p11_mult_21_n276), .CO(p11_mult_21_n271), .S(p11_mult_21_n272) );
  FA_X1 p11_mult_21_U122 ( .A(p11_mult_21_n281), .B(p11_mult_21_n283), .CI(
        p11_mult_21_n274), .CO(p11_mult_21_n269), .S(p11_mult_21_n270) );
  FA_X1 p11_mult_21_U121 ( .A(p11_mult_21_n279), .B(p11_mult_21_n272), .CI(
        p11_mult_21_n270), .CO(p11_mult_21_n267), .S(p11_mult_21_n268) );
  FA_X1 p11_mult_21_U120 ( .A(p11_mult_21_n361), .B(p11_mult_21_n337), .CI(
        p11_mult_21_n410), .CO(p11_mult_21_n265), .S(p11_mult_21_n266) );
  FA_X1 p11_mult_21_U109 ( .A(p11_mult_21_n349), .B(p11_mult_21_n397), .CI(
        p11_mult_21_n373), .CO(p11_mult_21_n263), .S(p11_mult_21_n264) );
  FA_X1 p11_mult_21_U108 ( .A(p11_mult_21_n275), .B(p11_mult_21_n385), .CI(
        p11_mult_21_n273), .CO(p11_mult_21_n261), .S(p11_mult_21_n262) );
  FA_X1 p11_mult_21_U107 ( .A(p11_mult_21_n264), .B(p11_mult_21_n266), .CI(
        p11_mult_21_n271), .CO(p11_mult_21_n259), .S(p11_mult_21_n260) );
  FA_X1 p11_mult_21_U106 ( .A(p11_mult_21_n262), .B(p11_mult_21_n269), .CI(
        p11_mult_21_n260), .CO(p11_mult_21_n257), .S(p11_mult_21_n258) );
  HA_X1 p11_mult_21_U105 ( .A(p11_mult_21_n317), .B(p11_mult_21_n336), .CO(
        p11_mult_21_n255), .S(p11_mult_21_n256) );
  FA_X1 p11_mult_21_U104 ( .A(p11_mult_21_n409), .B(p11_mult_21_n372), .CI(
        p11_mult_21_n396), .CO(p11_mult_21_n253), .S(p11_mult_21_n254) );
  FA_X1 p11_mult_21_U103 ( .A(p11_mult_21_n348), .B(p11_mult_21_n384), .CI(
        p11_mult_21_n360), .CO(p11_mult_21_n251), .S(p11_mult_21_n252) );
  FA_X1 p11_mult_21_U102 ( .A(p11_mult_21_n265), .B(p11_mult_21_n256), .CI(
        p11_mult_21_n263), .CO(p11_mult_21_n249), .S(p11_mult_21_n250) );
  FA_X1 p11_mult_21_U101 ( .A(p11_mult_21_n254), .B(p11_mult_21_n252), .CI(
        p11_mult_21_n261), .CO(p11_mult_21_n247), .S(p11_mult_21_n248) );
  FA_X1 p11_mult_21_U100 ( .A(p11_mult_21_n259), .B(p11_mult_21_n250), .CI(
        p11_mult_21_n248), .CO(p11_mult_21_n245), .S(p11_mult_21_n246) );
  FA_X1 p11_mult_21_U97 ( .A(p11_mult_21_n395), .B(p11_mult_21_n359), .CI(
        p11_mult_21_n408), .CO(p11_mult_21_n241), .S(p11_mult_21_n242) );
  FA_X1 p11_mult_21_U96 ( .A(p11_mult_21_n335), .B(p11_mult_21_n371), .CI(
        p11_mult_21_n255), .CO(p11_mult_21_n239), .S(p11_mult_21_n240) );
  FA_X1 p11_mult_21_U95 ( .A(p11_mult_21_n253), .B(p11_mult_21_n244), .CI(
        p11_mult_21_n251), .CO(p11_mult_21_n237), .S(p11_mult_21_n238) );
  FA_X1 p11_mult_21_U94 ( .A(p11_mult_21_n240), .B(p11_mult_21_n242), .CI(
        p11_mult_21_n249), .CO(p11_mult_21_n235), .S(p11_mult_21_n236) );
  FA_X1 p11_mult_21_U93 ( .A(p11_mult_21_n247), .B(p11_mult_21_n238), .CI(
        p11_mult_21_n236), .CO(p11_mult_21_n233), .S(p11_mult_21_n234) );
  FA_X1 p11_mult_21_U91 ( .A(p11_mult_21_n382), .B(p11_mult_21_n346), .CI(
        p11_mult_21_n232), .CO(p11_mult_21_n229), .S(p11_mult_21_n230) );
  FA_X1 p11_mult_21_U90 ( .A(p11_mult_21_n334), .B(p11_mult_21_n370), .CI(
        p11_mult_21_n358), .CO(p11_mult_21_n227), .S(p11_mult_21_n228) );
  FA_X1 p11_mult_21_U89 ( .A(p11_mult_21_n241), .B(p11_mult_21_n243), .CI(
        p11_mult_21_n239), .CO(p11_mult_21_n225), .S(p11_mult_21_n226) );
  FA_X1 p11_mult_21_U88 ( .A(p11_mult_21_n230), .B(p11_mult_21_n228), .CI(
        p11_mult_21_n237), .CO(p11_mult_21_n223), .S(p11_mult_21_n224) );
  FA_X1 p11_mult_21_U87 ( .A(p11_mult_21_n235), .B(p11_mult_21_n226), .CI(
        p11_mult_21_n224), .CO(p11_mult_21_n221), .S(p11_mult_21_n222) );
  FA_X1 p11_mult_21_U86 ( .A(p11_mult_21_n231), .B(p11_mult_21_n333), .CI(
        p11_mult_21_n394), .CO(p11_mult_21_n219), .S(p11_mult_21_n220) );
  FA_X1 p11_mult_21_U85 ( .A(p11_mult_21_n345), .B(p11_mult_21_n381), .CI(
        p11_mult_21_n357), .CO(p11_mult_21_n217), .S(p11_mult_21_n218) );
  FA_X1 p11_mult_21_U84 ( .A(p11_mult_21_n229), .B(p11_mult_21_n369), .CI(
        p11_mult_21_n227), .CO(p11_mult_21_n215), .S(p11_mult_21_n216) );
  FA_X1 p11_mult_21_U83 ( .A(p11_mult_21_n220), .B(p11_mult_21_n218), .CI(
        p11_mult_21_n225), .CO(p11_mult_21_n213), .S(p11_mult_21_n214) );
  FA_X1 p11_mult_21_U82 ( .A(p11_mult_21_n223), .B(p11_mult_21_n216), .CI(
        p11_mult_21_n214), .CO(p11_mult_21_n211), .S(p11_mult_21_n212) );
  FA_X1 p11_mult_21_U80 ( .A(p11_mult_21_n368), .B(p11_mult_21_n344), .CI(
        p11_mult_21_n210), .CO(p11_mult_21_n207), .S(p11_mult_21_n208) );
  FA_X1 p11_mult_21_U79 ( .A(p11_mult_21_n332), .B(p11_mult_21_n356), .CI(
        p11_mult_21_n219), .CO(p11_mult_21_n205), .S(p11_mult_21_n206) );
  FA_X1 p11_mult_21_U78 ( .A(p11_mult_21_n208), .B(p11_mult_21_n217), .CI(
        p11_mult_21_n215), .CO(p11_mult_21_n203), .S(p11_mult_21_n204) );
  FA_X1 p11_mult_21_U77 ( .A(p11_mult_21_n213), .B(p11_mult_21_n206), .CI(
        p11_mult_21_n204), .CO(p11_mult_21_n201), .S(p11_mult_21_n202) );
  FA_X1 p11_mult_21_U76 ( .A(p11_mult_21_n209), .B(p11_mult_21_n331), .CI(
        p11_mult_21_n380), .CO(p11_mult_21_n199), .S(p11_mult_21_n200) );
  FA_X1 p11_mult_21_U75 ( .A(p11_mult_21_n355), .B(p11_mult_21_n343), .CI(
        p11_mult_21_n367), .CO(p11_mult_21_n197), .S(p11_mult_21_n198) );
  FA_X1 p11_mult_21_U74 ( .A(p11_mult_21_n198), .B(p11_mult_21_n207), .CI(
        p11_mult_21_n200), .CO(p11_mult_21_n195), .S(p11_mult_21_n196) );
  FA_X1 p11_mult_21_U73 ( .A(p11_mult_21_n203), .B(p11_mult_21_n205), .CI(
        p11_mult_21_n196), .CO(p11_mult_21_n193), .S(p11_mult_21_n194) );
  FA_X1 p11_mult_21_U71 ( .A(p11_mult_21_n330), .B(p11_mult_21_n342), .CI(
        p11_mult_21_n192), .CO(p11_mult_21_n189), .S(p11_mult_21_n190) );
  FA_X1 p11_mult_21_U70 ( .A(p11_mult_21_n199), .B(p11_mult_21_n354), .CI(
        p11_mult_21_n197), .CO(p11_mult_21_n187), .S(p11_mult_21_n188) );
  FA_X1 p11_mult_21_U69 ( .A(p11_mult_21_n188), .B(p11_mult_21_n190), .CI(
        p11_mult_21_n195), .CO(p11_mult_21_n185), .S(p11_mult_21_n186) );
  FA_X1 p11_mult_21_U68 ( .A(p11_mult_21_n191), .B(p11_mult_21_n329), .CI(
        p11_mult_21_n366), .CO(p11_mult_21_n183), .S(p11_mult_21_n184) );
  FA_X1 p11_mult_21_U67 ( .A(p11_mult_21_n341), .B(p11_mult_21_n353), .CI(
        p11_mult_21_n189), .CO(p11_mult_21_n181), .S(p11_mult_21_n182) );
  FA_X1 p11_mult_21_U66 ( .A(p11_mult_21_n187), .B(p11_mult_21_n184), .CI(
        p11_mult_21_n182), .CO(p11_mult_21_n179), .S(p11_mult_21_n180) );
  FA_X1 p11_mult_21_U64 ( .A(p11_mult_21_n328), .B(p11_mult_21_n340), .CI(
        p11_mult_21_n178), .CO(p11_mult_21_n175), .S(p11_mult_21_n176) );
  FA_X1 p11_mult_21_U63 ( .A(p11_mult_21_n176), .B(p11_mult_21_n183), .CI(
        p11_mult_21_n181), .CO(p11_mult_21_n173), .S(p11_mult_21_n174) );
  FA_X1 p11_mult_21_U62 ( .A(p11_mult_21_n327), .B(p11_mult_21_n177), .CI(
        p11_mult_21_n352), .CO(p11_mult_21_n171), .S(p11_mult_21_n172) );
  FA_X1 p11_mult_21_U61 ( .A(p11_mult_21_n175), .B(p11_mult_21_n339), .CI(
        p11_mult_21_n172), .CO(p11_mult_21_n169), .S(p11_mult_21_n170) );
  FA_X1 p11_mult_21_U59 ( .A(p11_mult_21_n168), .B(p11_mult_21_n326), .CI(
        p11_mult_21_n171), .CO(p11_mult_21_n165), .S(p11_mult_21_n166) );
  FA_X1 p11_mult_21_U58 ( .A(p11_mult_21_n325), .B(p11_mult_21_n167), .CI(
        p11_mult_21_n338), .CO(p11_mult_21_n163), .S(p11_mult_21_n164) );
  FA_X1 p11_mult_21_U41 ( .A(p11_mult_21_n212), .B(p11_mult_21_n221), .CI(
        p11_mult_21_n146), .CO(p11_mult_21_n145), .S(temp6[3]) );
  FA_X1 p11_mult_21_U40 ( .A(p11_mult_21_n202), .B(p11_mult_21_n211), .CI(
        p11_mult_21_n145), .CO(p11_mult_21_n144), .S(temp6[4]) );
  FA_X1 p11_mult_21_U39 ( .A(p11_mult_21_n194), .B(p11_mult_21_n201), .CI(
        p11_mult_21_n144), .CO(p11_mult_21_n143), .S(temp6[5]) );
  FA_X1 p11_mult_21_U37 ( .A(p11_mult_21_n180), .B(p11_mult_21_n185), .CI(
        p11_mult_21_n142), .CO(p11_mult_21_n141), .S(temp6[7]) );
  FA_X1 p11_mult_21_U30 ( .A(p11_mult_21_n174), .B(p11_mult_21_n179), .CI(
        p11_mult_21_n141), .CO(p11_mult_21_n140), .S(temp6[8]) );
  FA_X1 p11_mult_21_U20 ( .A(p11_mult_21_n170), .B(p11_mult_21_n173), .CI(
        p11_mult_21_n140), .CO(p11_mult_21_n139), .S(temp6[9]) );
  FA_X1 p11_mult_21_U10 ( .A(p11_mult_21_n166), .B(p11_mult_21_n169), .CI(
        p11_mult_21_n139), .CO(p11_mult_21_n138), .S(temp6[10]) );
  FA_X1 p11_mult_21_U9 ( .A(p11_mult_21_n165), .B(p11_mult_21_n164), .CI(
        p11_mult_21_n138), .CO(p11_mult_21_n137), .S(temp6[11]) );
  FA_X1 p11_mult_21_U8 ( .A(p11_mult_21_n163), .B(p11_mult_21_n162), .CI(
        p11_mult_21_n137), .CO(p11_mult_21_n136), .S(temp6[12]) );
  INV_X1 p10_mult_21_U438 ( .A(p10_mult_21_n875), .ZN(p10_mult_21_n873) );
  INV_X1 p10_mult_21_U453 ( .A(p10_mult_21_n901), .ZN(p10_mult_21_n899) );
  INV_X1 p10_mult_21_U463 ( .A(p10_mult_21_n915), .ZN(p10_mult_21_n914) );
  INV_X1 p10_mult_21_U484 ( .A(p10_mult_21_n947), .ZN(p10_mult_21_n945) );
  INV_X1 p10_mult_21_U494 ( .A(p10_mult_21_n963), .ZN(p10_mult_21_n962) );
  INV_X1 p10_mult_21_U496 ( .A(p10_mult_21_n966), .ZN(p10_mult_21_n965) );
  INV_X1 p10_mult_21_U562 ( .A(p10_mult_21_n1059), .ZN(p10_mult_21_n1058) );
  INV_X1 p10_mult_21_U566 ( .A(p10_mult_21_n1061), .ZN(p10_mult_21_n1060) );
  INV_X1 p10_mult_21_U652 ( .A(p10_mult_21_n1194), .ZN(p10_mult_21_n1191) );
  INV_X1 p10_mult_21_U661 ( .A(p10_mult_21_n1219), .ZN(p10_mult_21_n1218) );
  INV_X1 p10_mult_21_U410 ( .A(p10_mult_21_n1243), .ZN(p10_mult_21_n837) );
  INV_X1 p10_mult_21_U709 ( .A(p10_mult_21_n1300), .ZN(p10_mult_21_n1299) );
  INV_X1 p10_mult_21_U418 ( .A(p10_mult_21_n1303), .ZN(p10_mult_21_n845) );
  INV_X1 p10_mult_21_U412 ( .A(p10_mult_21_n1271), .ZN(p10_mult_21_n839) );
  INV_X1 p10_mult_21_U414 ( .A(p10_mult_21_n1286), .ZN(p10_mult_21_n841) );
  INV_X1 p10_mult_21_U726 ( .A(p10_mult_21_n1309), .ZN(p10_mult_21_n1209) );
  INV_X1 p10_mult_21_U422 ( .A(p10_mult_21_n1310), .ZN(p10_mult_21_n849) );
  INV_X1 p10_mult_21_U745 ( .A(p10_mult_21_n985), .ZN(p10_mult_21_n952) );
  INV_X1 p10_mult_21_U750 ( .A(p10_mult_21_n1330), .ZN(p10_mult_21_n1201) );
  INV_X1 p10_mult_21_U837 ( .A(p10_mult_21_n1352), .ZN(p10_mult_21_n1387) );
  INV_X1 p10_mult_21_U785 ( .A(p10_mult_21_n1362), .ZN(p10_mult_21_n1356) );
  INV_X1 p10_mult_21_U835 ( .A(p10_mult_21_n1386), .ZN(p10_mult_21_n1383) );
  INV_X1 p10_mult_21_U578 ( .A(p10_mult_21_n1084), .ZN(p10_mult_21_n1083) );
  INV_X1 p10_mult_21_U581 ( .A(p10_mult_21_n1086), .ZN(p10_mult_21_n1085) );
  INV_X1 p10_mult_21_U705 ( .A(p10_mult_21_n1113), .ZN(p10_mult_21_n1090) );
  AND2_X1 p10_mult_21_U611 ( .A1(p10_mult_21_n1123), .A2(p10_mult_21_n1124), 
        .ZN(p10_mult_21_n1097) );
  AND2_X1 p10_mult_21_U640 ( .A1(p10_mult_21_n1172), .A2(p10_mult_21_n1173), 
        .ZN(p10_mult_21_n1128) );
  INV_X1 p10_mult_21_U868 ( .A(A2[1]), .ZN(p10_mult_21_n1298) );
  INV_X1 p10_mult_21_U571 ( .A(p10_mult_21_n1070), .ZN(p10_mult_21_n1052) );
  INV_X1 p10_mult_21_U630 ( .A(p10_mult_21_n1158), .ZN(p10_mult_21_n1157) );
  INV_X1 p10_mult_21_U881 ( .A(A2[4]), .ZN(p10_mult_21_n1094) );
  INV_X1 p10_mult_21_U801 ( .A(p10_mult_21_n1360), .ZN(p10_mult_21_n1369) );
  INV_X1 p10_mult_21_U872 ( .A(A2[2]), .ZN(p10_mult_21_n1175) );
  INV_X1 p10_mult_21_U869 ( .A(p10_mult_21_n903), .ZN(p10_mult_21_n881) );
  INV_X1 p10_mult_21_U873 ( .A(p10_mult_21_n911), .ZN(p10_mult_21_n880) );
  INV_X1 p10_mult_21_U627 ( .A(p10_mult_21_n1151), .ZN(p10_mult_21_n1107) );
  INV_X1 p10_mult_21_U814 ( .A(p10_mult_21_n1167), .ZN(p10_mult_21_n1373) );
  INV_X1 p10_mult_21_U744 ( .A(p10_mult_21_n1014), .ZN(p10_mult_21_n951) );
  INV_X1 p10_mult_21_U519 ( .A(p10_mult_21_n994), .ZN(p10_mult_21_n992) );
  INV_X1 p10_mult_21_U521 ( .A(p10_mult_21_n998), .ZN(p10_mult_21_n995) );
  INV_X1 p10_mult_21_U850 ( .A(A2[5]), .ZN(p10_mult_21_n1062) );
  INV_X1 p10_mult_21_U827 ( .A(p10_mult_21_n1092), .ZN(p10_mult_21_n863) );
  INV_X1 p10_mult_21_U568 ( .A(p10_mult_21_n1063), .ZN(p10_mult_21_n862) );
  INV_X1 p10_mult_21_U843 ( .A(A2[8]), .ZN(p10_mult_21_n955) );
  INV_X1 p10_mult_21_U859 ( .A(A2[9]), .ZN(p10_mult_21_n935) );
  INV_X1 p10_mult_21_U766 ( .A(p10_mult_21_n937), .ZN(p10_mult_21_n918) );
  INV_X1 p10_mult_21_U765 ( .A(p10_mult_21_n964), .ZN(p10_mult_21_n917) );
  INV_X1 p10_mult_21_U533 ( .A(p10_mult_21_n1016), .ZN(p10_mult_21_n999) );
  INV_X1 p10_mult_21_U535 ( .A(p10_mult_21_n993), .ZN(p10_mult_21_n1019) );
  INV_X1 p10_mult_21_U816 ( .A(A2[13]), .ZN(p10_mult_21_n868) );
  INV_X1 p10_mult_21_U894 ( .A(A2[12]), .ZN(p10_mult_21_n879) );
  INV_X1 p10_mult_21_U853 ( .A(A2[6]), .ZN(p10_mult_21_n1025) );
  INV_X1 p10_mult_21_U819 ( .A(A2[7]), .ZN(p10_mult_21_n983) );
  INV_X1 p10_mult_21_U863 ( .A(A2[10]), .ZN(p10_mult_21_n921) );
  INV_X1 p10_mult_21_U822 ( .A(A2[11]), .ZN(p10_mult_21_n897) );
  OAI22_X1 p10_mult_21_U874 ( .A1(n901), .A2(n912), .B1(reg4[10]), .B2(reg4[9]), .ZN(p10_mult_21_n911) );
  OAI22_X1 p10_mult_21_U883 ( .A1(n908), .A2(n904), .B1(reg4[7]), .B2(reg4[8]), 
        .ZN(p10_mult_21_n964) );
  XNOR2_X1 p10_mult_21_U620 ( .A(p10_mult_21_n1137), .B(p10_mult_21_n1139), 
        .ZN(p10_mult_21_n1140) );
  XNOR2_X1 p10_mult_21_U645 ( .A(p10_mult_21_n1143), .B(p10_mult_21_n1177), 
        .ZN(temp5[0]) );
  XNOR2_X1 p10_mult_21_U570 ( .A(p10_mult_21_n1067), .B(p10_mult_21_n1035), 
        .ZN(temp5[3]) );
  XNOR2_X1 p10_mult_21_U543 ( .A(p10_mult_21_n1028), .B(p10_mult_21_n1032), 
        .ZN(temp5[4]) );
  XNOR2_X1 p10_mult_21_U523 ( .A(p10_mult_21_n1002), .B(p10_mult_21_n976), 
        .ZN(temp5[5]) );
  XNOR2_X1 p10_mult_21_U501 ( .A(p10_mult_21_n969), .B(p10_mult_21_n973), .ZN(
        temp5[6]) );
  XNOR2_X1 p10_mult_21_U485 ( .A(p10_mult_21_n948), .B(p10_mult_21_n928), .ZN(
        temp5[7]) );
  XNOR2_X1 p10_mult_21_U459 ( .A(p10_mult_21_n889), .B(p10_mult_21_n890), .ZN(
        p10_mult_21_n906) );
  XNOR2_X1 p10_mult_21_U469 ( .A(p10_mult_21_n909), .B(p10_mult_21_n925), .ZN(
        temp5[8]) );
  XNOR2_X1 p10_mult_21_U447 ( .A(p10_mult_21_n885), .B(p10_mult_21_n888), .ZN(
        temp5[10]) );
  AOI222_X1 p10_mult_21_U437 ( .A1(p10_mult_21_n872), .A2(p10_mult_21_n873), 
        .B1(p10_mult_21_n872), .B2(p10_mult_21_n874), .C1(p10_mult_21_n873), 
        .C2(p10_mult_21_n874), .ZN(p10_mult_21_n857) );
  AOI22_X1 p10_mult_21_U433 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n864), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n866), .ZN(p10_mult_21_n860) );
  AOI22_X1 p10_mult_21_U434 ( .A1(A2[13]), .A2(reg4[13]), .B1(n903), .B2(
        p10_mult_21_n868), .ZN(p10_mult_21_n864) );
  XNOR2_X1 p10_mult_21_U440 ( .A(p10_mult_21_n874), .B(p10_mult_21_n875), .ZN(
        p10_mult_21_n877) );
  AOI22_X1 p10_mult_21_U441 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n866), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n878), .ZN(p10_mult_21_n875) );
  OAI22_X1 p10_mult_21_U442 ( .A1(n903), .A2(A2[12]), .B1(p10_mult_21_n879), 
        .B2(reg4[13]), .ZN(p10_mult_21_n866) );
  OAI21_X1 p10_mult_21_U443 ( .B1(p10_mult_21_n880), .B2(p10_mult_21_n881), 
        .A(p10_mult_21_n882), .ZN(p10_mult_21_n872) );
  AOI222_X1 p10_mult_21_U446 ( .A1(p10_mult_21_n886), .A2(p10_mult_21_n887), 
        .B1(p10_mult_21_n886), .B2(p10_mult_21_n874), .C1(p10_mult_21_n887), 
        .C2(p10_mult_21_n874), .ZN(p10_mult_21_n869) );
  AOI22_X1 p10_mult_21_U450 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n878), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n896), .ZN(p10_mult_21_n887) );
  OAI22_X1 p10_mult_21_U451 ( .A1(n903), .A2(A2[11]), .B1(p10_mult_21_n897), 
        .B2(reg4[13]), .ZN(p10_mult_21_n878) );
  AOI222_X1 p10_mult_21_U452 ( .A1(p10_mult_21_n898), .A2(p10_mult_21_n899), 
        .B1(p10_mult_21_n898), .B2(p10_mult_21_n900), .C1(p10_mult_21_n899), 
        .C2(p10_mult_21_n900), .ZN(p10_mult_21_n886) );
  OAI21_X1 p10_mult_21_U454 ( .B1(p10_mult_21_n902), .B2(p10_mult_21_n903), 
        .A(p10_mult_21_n904), .ZN(p10_mult_21_n874) );
  NAND2_X1 p10_mult_21_U455 ( .A1(p10_mult_21_n880), .A2(p10_mult_21_n882), 
        .ZN(p10_mult_21_n904) );
  AOI22_X1 p10_mult_21_U456 ( .A1(A2[13]), .A2(reg4[11]), .B1(n902), .B2(
        p10_mult_21_n868), .ZN(p10_mult_21_n882) );
  AOI222_X1 p10_mult_21_U449 ( .A1(p10_mult_21_n892), .A2(p10_mult_21_n893), 
        .B1(p10_mult_21_n892), .B2(p10_mult_21_n894), .C1(p10_mult_21_n893), 
        .C2(p10_mult_21_n894), .ZN(p10_mult_21_n883) );
  OAI22_X1 p10_mult_21_U460 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n902), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n912), .ZN(p10_mult_21_n893) );
  AOI22_X1 p10_mult_21_U461 ( .A1(reg4[11]), .A2(p10_mult_21_n879), .B1(A2[12]), .B2(n902), .ZN(p10_mult_21_n902) );
  AOI222_X1 p10_mult_21_U462 ( .A1(p10_mult_21_n913), .A2(p10_mult_21_n914), 
        .B1(p10_mult_21_n913), .B2(p10_mult_21_n900), .C1(p10_mult_21_n914), 
        .C2(p10_mult_21_n900), .ZN(p10_mult_21_n892) );
  OAI21_X1 p10_mult_21_U464 ( .B1(p10_mult_21_n917), .B2(p10_mult_21_n918), 
        .A(p10_mult_21_n919), .ZN(p10_mult_21_n898) );
  XNOR2_X1 p10_mult_21_U465 ( .A(p10_mult_21_n900), .B(p10_mult_21_n901), .ZN(
        p10_mult_21_n916) );
  AOI22_X1 p10_mult_21_U466 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n896), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n920), .ZN(p10_mult_21_n901) );
  OAI22_X1 p10_mult_21_U467 ( .A1(n903), .A2(A2[10]), .B1(p10_mult_21_n921), 
        .B2(reg4[13]), .ZN(p10_mult_21_n896) );
  AOI222_X1 p10_mult_21_U471 ( .A1(p10_mult_21_n929), .A2(p10_mult_21_n930), 
        .B1(p10_mult_21_n929), .B2(p10_mult_21_n931), .C1(p10_mult_21_n930), 
        .C2(p10_mult_21_n931), .ZN(p10_mult_21_n907) );
  XNOR2_X1 p10_mult_21_U472 ( .A(p10_mult_21_n932), .B(p10_mult_21_n924), .ZN(
        p10_mult_21_n909) );
  XNOR2_X1 p10_mult_21_U473 ( .A(p10_mult_21_n915), .B(p10_mult_21_n933), .ZN(
        p10_mult_21_n924) );
  AOI22_X1 p10_mult_21_U474 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n920), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n934), .ZN(p10_mult_21_n913) );
  OAI22_X1 p10_mult_21_U475 ( .A1(n903), .A2(A2[9]), .B1(p10_mult_21_n935), 
        .B2(reg4[13]), .ZN(p10_mult_21_n920) );
  OAI21_X1 p10_mult_21_U476 ( .B1(p10_mult_21_n936), .B2(p10_mult_21_n937), 
        .A(p10_mult_21_n938), .ZN(p10_mult_21_n900) );
  NAND2_X1 p10_mult_21_U477 ( .A1(p10_mult_21_n917), .A2(p10_mult_21_n919), 
        .ZN(p10_mult_21_n938) );
  AOI22_X1 p10_mult_21_U478 ( .A1(A2[13]), .A2(reg4[9]), .B1(n901), .B2(
        p10_mult_21_n868), .ZN(p10_mult_21_n919) );
  OAI22_X1 p10_mult_21_U479 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n912), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n940), .ZN(p10_mult_21_n915) );
  OAI22_X1 p10_mult_21_U480 ( .A1(n902), .A2(p10_mult_21_n897), .B1(A2[11]), 
        .B2(reg4[11]), .ZN(p10_mult_21_n912) );
  XNOR2_X1 p10_mult_21_U481 ( .A(p10_mult_21_n922), .B(p10_mult_21_n923), .ZN(
        p10_mult_21_n932) );
  AOI222_X1 p10_mult_21_U482 ( .A1(p10_mult_21_n941), .A2(p10_mult_21_n942), 
        .B1(p10_mult_21_n941), .B2(p10_mult_21_n943), .C1(p10_mult_21_n942), 
        .C2(p10_mult_21_n943), .ZN(p10_mult_21_n923) );
  AOI222_X1 p10_mult_21_U483 ( .A1(p10_mult_21_n944), .A2(p10_mult_21_n945), 
        .B1(p10_mult_21_n944), .B2(p10_mult_21_n946), .C1(p10_mult_21_n945), 
        .C2(p10_mult_21_n946), .ZN(p10_mult_21_n922) );
  OAI21_X1 p10_mult_21_U486 ( .B1(p10_mult_21_n951), .B2(p10_mult_21_n952), 
        .A(p10_mult_21_n953), .ZN(p10_mult_21_n944) );
  XNOR2_X1 p10_mult_21_U487 ( .A(p10_mult_21_n946), .B(p10_mult_21_n947), .ZN(
        p10_mult_21_n950) );
  AOI22_X1 p10_mult_21_U488 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n934), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n954), .ZN(p10_mult_21_n947) );
  AOI22_X1 p10_mult_21_U489 ( .A1(reg4[13]), .A2(A2[8]), .B1(p10_mult_21_n955), 
        .B2(n903), .ZN(p10_mult_21_n934) );
  AOI222_X1 p10_mult_21_U490 ( .A1(p10_mult_21_n956), .A2(p10_mult_21_n957), 
        .B1(p10_mult_21_n956), .B2(p10_mult_21_n958), .C1(p10_mult_21_n957), 
        .C2(p10_mult_21_n958), .ZN(p10_mult_21_n929) );
  OAI22_X1 p10_mult_21_U491 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n940), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n960), .ZN(p10_mult_21_n942) );
  OAI22_X1 p10_mult_21_U492 ( .A1(n902), .A2(p10_mult_21_n921), .B1(A2[10]), 
        .B2(reg4[11]), .ZN(p10_mult_21_n940) );
  AOI222_X1 p10_mult_21_U493 ( .A1(p10_mult_21_n961), .A2(p10_mult_21_n962), 
        .B1(p10_mult_21_n961), .B2(p10_mult_21_n946), .C1(p10_mult_21_n962), 
        .C2(p10_mult_21_n946), .ZN(p10_mult_21_n941) );
  OAI22_X1 p10_mult_21_U495 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n936), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n965), .ZN(p10_mult_21_n943) );
  AOI22_X1 p10_mult_21_U497 ( .A1(A2[12]), .A2(n901), .B1(reg4[9]), .B2(
        p10_mult_21_n879), .ZN(p10_mult_21_n936) );
  XNOR2_X1 p10_mult_21_U513 ( .A(p10_mult_21_n970), .B(p10_mult_21_n971), .ZN(
        p10_mult_21_n980) );
  AOI222_X1 p10_mult_21_U524 ( .A1(p10_mult_21_n1004), .A2(p10_mult_21_n1005), 
        .B1(p10_mult_21_n1004), .B2(p10_mult_21_n1006), .C1(p10_mult_21_n1005), 
        .C2(p10_mult_21_n1006), .ZN(p10_mult_21_n978) );
  AOI222_X1 p10_mult_21_U525 ( .A1(p10_mult_21_n1007), .A2(p10_mult_21_n1008), 
        .B1(p10_mult_21_n1007), .B2(p10_mult_21_n1009), .C1(p10_mult_21_n1008), 
        .C2(p10_mult_21_n1009), .ZN(p10_mult_21_n977) );
  AOI222_X1 p10_mult_21_U542 ( .A1(p10_mult_21_n1029), .A2(p10_mult_21_n1030), 
        .B1(p10_mult_21_n1029), .B2(p10_mult_21_n1031), .C1(p10_mult_21_n1030), 
        .C2(p10_mult_21_n1031), .ZN(p10_mult_21_n974) );
  XNOR2_X1 p10_mult_21_U546 ( .A(p10_mult_21_n1040), .B(p10_mult_21_n1006), 
        .ZN(p10_mult_21_n1031) );
  XNOR2_X1 p10_mult_21_U547 ( .A(p10_mult_21_n1018), .B(p10_mult_21_n1041), 
        .ZN(p10_mult_21_n1006) );
  XNOR2_X1 p10_mult_21_U548 ( .A(p10_mult_21_n993), .B(p10_mult_21_n1017), 
        .ZN(p10_mult_21_n1041) );
  XNOR2_X1 p10_mult_21_U556 ( .A(p10_mult_21_n1004), .B(p10_mult_21_n1005), 
        .ZN(p10_mult_21_n1040) );
  AOI222_X1 p10_mult_21_U557 ( .A1(p10_mult_21_n1048), .A2(p10_mult_21_n1049), 
        .B1(p10_mult_21_n1048), .B2(p10_mult_21_n1050), .C1(p10_mult_21_n1049), 
        .C2(p10_mult_21_n1050), .ZN(p10_mult_21_n1005) );
  AOI222_X1 p10_mult_21_U558 ( .A1(p10_mult_21_n1051), .A2(p10_mult_21_n1052), 
        .B1(p10_mult_21_n1051), .B2(p10_mult_21_n1053), .C1(p10_mult_21_n1052), 
        .C2(p10_mult_21_n1053), .ZN(p10_mult_21_n1004) );
  AOI222_X1 p10_mult_21_U559 ( .A1(p10_mult_21_n1054), .A2(p10_mult_21_n1055), 
        .B1(p10_mult_21_n1054), .B2(p10_mult_21_n1056), .C1(p10_mult_21_n1055), 
        .C2(p10_mult_21_n1056), .ZN(p10_mult_21_n1029) );
  XNOR2_X1 p10_mult_21_U560 ( .A(p10_mult_21_n1057), .B(p10_mult_21_n1009), 
        .ZN(p10_mult_21_n1030) );
  AOI22_X1 p10_mult_21_U561 ( .A1(p10_mult_21_n917), .A2(p10_mult_21_n1013), 
        .B1(p10_mult_21_n918), .B2(p10_mult_21_n1058), .ZN(p10_mult_21_n1009)
         );
  XNOR2_X1 p10_mult_21_U564 ( .A(p10_mult_21_n1007), .B(p10_mult_21_n1008), 
        .ZN(p10_mult_21_n1057) );
  AOI22_X1 p10_mult_21_U565 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n1024), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n1060), .ZN(p10_mult_21_n1008)
         );
  AOI222_X1 p10_mult_21_U569 ( .A1(p10_mult_21_n1064), .A2(p10_mult_21_n1065), 
        .B1(p10_mult_21_n1064), .B2(p10_mult_21_n1066), .C1(p10_mult_21_n1065), 
        .C2(p10_mult_21_n1066), .ZN(p10_mult_21_n1007) );
  AOI222_X1 p10_mult_21_U621 ( .A1(p10_mult_21_n1144), .A2(p10_mult_21_n1145), 
        .B1(p10_mult_21_n1144), .B2(p10_mult_21_n1146), .C1(p10_mult_21_n1145), 
        .C2(p10_mult_21_n1146), .ZN(p10_mult_21_n1139) );
  AOI222_X1 p10_mult_21_U651 ( .A1(p10_mult_21_n1191), .A2(p10_mult_21_n1192), 
        .B1(p10_mult_21_n1191), .B2(p10_mult_21_n1193), .C1(p10_mult_21_n1192), 
        .C2(p10_mult_21_n1193), .ZN(p10_mult_21_n1190) );
  XNOR2_X1 p10_mult_21_U654 ( .A(p10_mult_21_n1198), .B(p10_mult_21_n1193), 
        .ZN(p10_mult_21_n1197) );
  XNOR2_X1 p10_mult_21_U655 ( .A(p10_mult_21_n1203), .B(p10_mult_21_n1204), 
        .ZN(p10_mult_21_n1192) );
  XNOR2_X1 p10_mult_21_U656 ( .A(p10_mult_21_n1205), .B(p10_mult_21_n1206), 
        .ZN(p10_mult_21_n1203) );
  AOI222_X1 p10_mult_21_U657 ( .A1(p10_mult_21_n1207), .A2(p10_mult_21_n1208), 
        .B1(p10_mult_21_n1207), .B2(p10_mult_21_n1209), .C1(p10_mult_21_n1208), 
        .C2(p10_mult_21_n1209), .ZN(p10_mult_21_n1194) );
  AOI222_X1 p10_mult_21_U658 ( .A1(p10_mult_21_n1210), .A2(p10_mult_21_n1211), 
        .B1(p10_mult_21_n1210), .B2(p10_mult_21_n1212), .C1(p10_mult_21_n1211), 
        .C2(p10_mult_21_n1212), .ZN(p10_mult_21_n1196) );
  AOI222_X1 p10_mult_21_U660 ( .A1(p10_mult_21_n1216), .A2(p10_mult_21_n1217), 
        .B1(p10_mult_21_n1216), .B2(p10_mult_21_n1218), .C1(p10_mult_21_n1217), 
        .C2(p10_mult_21_n1218), .ZN(p10_mult_21_n1215) );
  XNOR2_X1 p10_mult_21_U663 ( .A(p10_mult_21_n1224), .B(p10_mult_21_n1225), 
        .ZN(p10_mult_21_n1217) );
  XNOR2_X1 p10_mult_21_U664 ( .A(p10_mult_21_n1226), .B(p10_mult_21_n1227), 
        .ZN(p10_mult_21_n1224) );
  AOI222_X1 p10_mult_21_U666 ( .A1(p10_mult_21_n1232), .A2(p10_mult_21_n1233), 
        .B1(p10_mult_21_n1232), .B2(p10_mult_21_n1234), .C1(p10_mult_21_n1233), 
        .C2(p10_mult_21_n1234), .ZN(p10_mult_21_n1219) );
  AOI222_X1 p10_mult_21_U667 ( .A1(p10_mult_21_n1235), .A2(p10_mult_21_n1236), 
        .B1(p10_mult_21_n1235), .B2(p10_mult_21_n1237), .C1(p10_mult_21_n1236), 
        .C2(p10_mult_21_n1237), .ZN(p10_mult_21_n1221) );
  XNOR2_X1 p10_mult_21_U670 ( .A(p10_mult_21_n1232), .B(p10_mult_21_n1234), 
        .ZN(p10_mult_21_n1242) );
  OAI22_X1 p10_mult_21_U671 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1246), 
        .B1(n735), .B2(p10_mult_21_n1247), .ZN(p10_mult_21_n1234) );
  AOI222_X1 p10_mult_21_U674 ( .A1(p10_mult_21_n1252), .A2(p10_mult_21_n1253), 
        .B1(p10_mult_21_n1252), .B2(p10_mult_21_n1254), .C1(p10_mult_21_n1253), 
        .C2(p10_mult_21_n1254), .ZN(p10_mult_21_n1235) );
  OAI22_X1 p10_mult_21_U708 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1247), 
        .B1(n735), .B2(p10_mult_21_n1299), .ZN(p10_mult_21_n1260) );
  AOI22_X1 p10_mult_21_U710 ( .A1(reg4[5]), .A2(p10_mult_21_n1175), .B1(A2[2]), 
        .B2(p10_mult_21_n1046), .ZN(p10_mult_21_n1247) );
  XNOR2_X1 p10_mult_21_U716 ( .A(p10_mult_21_n1302), .B(p10_mult_21_n1254), 
        .ZN(p10_mult_21_n1258) );
  XNOR2_X1 p10_mult_21_U718 ( .A(p10_mult_21_n1253), .B(p10_mult_21_n1252), 
        .ZN(p10_mult_21_n1302) );
  OAI22_X1 p10_mult_21_U697 ( .A1(A2[1]), .A2(p10_mult_21_n1294), .B1(
        p10_mult_21_n1295), .B2(n906), .ZN(p10_mult_21_n1293) );
  XNOR2_X1 p10_mult_21_U723 ( .A(p10_mult_21_n1304), .B(p10_mult_21_n1212), 
        .ZN(p10_mult_21_n1213) );
  XNOR2_X1 p10_mult_21_U724 ( .A(p10_mult_21_n1305), .B(p10_mult_21_n1208), 
        .ZN(p10_mult_21_n1212) );
  AOI222_X1 p10_mult_21_U727 ( .A1(p10_mult_21_n1227), .A2(p10_mult_21_n1226), 
        .B1(p10_mult_21_n1227), .B2(p10_mult_21_n1225), .C1(p10_mult_21_n1226), 
        .C2(p10_mult_21_n1225), .ZN(p10_mult_21_n1309) );
  OAI22_X1 p10_mult_21_U729 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1311), 
        .B1(n735), .B2(p10_mult_21_n1246), .ZN(p10_mult_21_n1226) );
  XNOR2_X1 p10_mult_21_U732 ( .A(p10_mult_21_n1211), .B(p10_mult_21_n1210), 
        .ZN(p10_mult_21_n1304) );
  XNOR2_X1 p10_mult_21_U733 ( .A(p10_mult_21_n1314), .B(p10_mult_21_n1315), 
        .ZN(p10_mult_21_n1312) );
  AOI222_X1 p10_mult_21_U734 ( .A1(p10_mult_21_n1231), .A2(p10_mult_21_n1230), 
        .B1(p10_mult_21_n1231), .B2(p10_mult_21_n1228), .C1(p10_mult_21_n1230), 
        .C2(p10_mult_21_n1228), .ZN(p10_mult_21_n1211) );
  OAI22_X1 p10_mult_21_U737 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1317), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1318), .ZN(p10_mult_21_n1230)
         );
  NOR2_X1 p10_mult_21_U738 ( .A1(p10_mult_21_n1251), .A2(p10_mult_21_n1250), 
        .ZN(p10_mult_21_n1231) );
  OAI22_X1 p10_mult_21_U742 ( .A1(n904), .A2(p10_mult_21_n1298), .B1(A2[1]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1318) );
  AOI222_X1 p10_mult_21_U649 ( .A1(p10_mult_21_n1185), .A2(p10_mult_21_n1186), 
        .B1(p10_mult_21_n1185), .B2(p10_mult_21_n1187), .C1(p10_mult_21_n1186), 
        .C2(p10_mult_21_n1187), .ZN(p10_mult_21_n1179) );
  XNOR2_X1 p10_mult_21_U748 ( .A(p10_mult_21_n1328), .B(p10_mult_21_n1329), 
        .ZN(p10_mult_21_n1326) );
  XNOR2_X1 p10_mult_21_U746 ( .A(p10_mult_21_n1322), .B(p10_mult_21_n1323), 
        .ZN(p10_mult_21_n1186) );
  XNOR2_X1 p10_mult_21_U747 ( .A(p10_mult_21_n1324), .B(p10_mult_21_n1325), 
        .ZN(p10_mult_21_n1322) );
  AOI222_X1 p10_mult_21_U749 ( .A1(p10_mult_21_n1199), .A2(p10_mult_21_n1202), 
        .B1(p10_mult_21_n1199), .B2(p10_mult_21_n1201), .C1(p10_mult_21_n1202), 
        .C2(p10_mult_21_n1201), .ZN(p10_mult_21_n1185) );
  OAI222_X1 p10_mult_21_U751 ( .A1(p10_mult_21_n1314), .A2(p10_mult_21_n1315), 
        .B1(p10_mult_21_n1314), .B2(p10_mult_21_n1313), .C1(p10_mult_21_n1315), 
        .C2(p10_mult_21_n1313), .ZN(p10_mult_21_n1330) );
  OAI22_X1 p10_mult_21_U754 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1332), 
        .B1(n735), .B2(p10_mult_21_n1311), .ZN(p10_mult_21_n1315) );
  OAI22_X1 p10_mult_21_U755 ( .A1(p10_mult_21_n1046), .A2(p10_mult_21_n1094), 
        .B1(A2[4]), .B2(reg4[5]), .ZN(p10_mult_21_n1311) );
  OAI22_X1 p10_mult_21_U756 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1333), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1317), .ZN(p10_mult_21_n1314)
         );
  OAI22_X1 p10_mult_21_U757 ( .A1(n904), .A2(p10_mult_21_n1175), .B1(A2[2]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1317) );
  XNOR2_X1 p10_mult_21_U758 ( .A(p10_mult_21_n1334), .B(p10_mult_21_n1335), 
        .ZN(p10_mult_21_n1202) );
  XNOR2_X1 p10_mult_21_U759 ( .A(p10_mult_21_n1336), .B(p10_mult_21_n1337), 
        .ZN(p10_mult_21_n1334) );
  NOR2_X1 p10_mult_21_U760 ( .A1(p10_mult_21_n1308), .A2(p10_mult_21_n1307), 
        .ZN(p10_mult_21_n1199) );
  XNOR2_X1 p10_mult_21_U647 ( .A(p10_mult_21_n1181), .B(p10_mult_21_n1182), 
        .ZN(p10_mult_21_n1180) );
  XNOR2_X1 p10_mult_21_U648 ( .A(p10_mult_21_n1183), .B(p10_mult_21_n1184), 
        .ZN(p10_mult_21_n1181) );
  AOI222_X1 p10_mult_21_U767 ( .A1(p10_mult_21_n1183), .A2(p10_mult_21_n1184), 
        .B1(p10_mult_21_n1183), .B2(p10_mult_21_n1182), .C1(p10_mult_21_n1184), 
        .C2(p10_mult_21_n1182), .ZN(p10_mult_21_n1142) );
  AOI222_X1 p10_mult_21_U768 ( .A1(p10_mult_21_n1324), .A2(p10_mult_21_n1325), 
        .B1(p10_mult_21_n1324), .B2(p10_mult_21_n1323), .C1(p10_mult_21_n1325), 
        .C2(p10_mult_21_n1323), .ZN(p10_mult_21_n1182) );
  XNOR2_X1 p10_mult_21_U769 ( .A(p10_mult_21_n1343), .B(p10_mult_21_n1344), 
        .ZN(p10_mult_21_n1341) );
  AOI222_X1 p10_mult_21_U770 ( .A1(p10_mult_21_n1337), .A2(p10_mult_21_n1336), 
        .B1(p10_mult_21_n1337), .B2(p10_mult_21_n1335), .C1(p10_mult_21_n1336), 
        .C2(p10_mult_21_n1335), .ZN(p10_mult_21_n1325) );
  OAI22_X1 p10_mult_21_U771 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1346), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1333), .ZN(p10_mult_21_n1336)
         );
  AOI222_X1 p10_mult_21_U774 ( .A1(p10_mult_21_n1205), .A2(p10_mult_21_n1206), 
        .B1(p10_mult_21_n1205), .B2(p10_mult_21_n1204), .C1(p10_mult_21_n1206), 
        .C2(p10_mult_21_n1204), .ZN(p10_mult_21_n1324) );
  OAI22_X1 p10_mult_21_U775 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1347), 
        .B1(n735), .B2(p10_mult_21_n1332), .ZN(p10_mult_21_n1204) );
  OAI22_X1 p10_mult_21_U776 ( .A1(p10_mult_21_n1046), .A2(p10_mult_21_n1062), 
        .B1(A2[5]), .B2(reg4[5]), .ZN(p10_mult_21_n1332) );
  OAI22_X1 p10_mult_21_U779 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1349), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1340), .ZN(p10_mult_21_n1205)
         );
  OAI22_X1 p10_mult_21_U780 ( .A1(n901), .A2(p10_mult_21_n1298), .B1(A2[1]), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1340) );
  XNOR2_X1 p10_mult_21_U781 ( .A(p10_mult_21_n1350), .B(p10_mult_21_n1351), 
        .ZN(p10_mult_21_n1184) );
  XNOR2_X1 p10_mult_21_U782 ( .A(p10_mult_21_n1359), .B(p10_mult_21_n1159), 
        .ZN(p10_mult_21_n1145) );
  XNOR2_X1 p10_mult_21_U796 ( .A(p10_mult_21_n1160), .B(p10_mult_21_n1161), 
        .ZN(p10_mult_21_n1359) );
  XNOR2_X1 p10_mult_21_U823 ( .A(p10_mult_21_n1377), .B(p10_mult_21_n1170), 
        .ZN(p10_mult_21_n1146) );
  XNOR2_X1 p10_mult_21_U832 ( .A(p10_mult_21_n1169), .B(p10_mult_21_n1168), 
        .ZN(p10_mult_21_n1377) );
  AOI222_X1 p10_mult_21_U836 ( .A1(p10_mult_21_n1351), .A2(p10_mult_21_n1353), 
        .B1(p10_mult_21_n1351), .B2(p10_mult_21_n1387), .C1(p10_mult_21_n1353), 
        .C2(p10_mult_21_n1387), .ZN(p10_mult_21_n1144) );
  AOI222_X1 p10_mult_21_U838 ( .A1(p10_mult_21_n1327), .A2(p10_mult_21_n1329), 
        .B1(p10_mult_21_n1327), .B2(p10_mult_21_n1328), .C1(p10_mult_21_n1329), 
        .C2(p10_mult_21_n1328), .ZN(p10_mult_21_n1352) );
  OAI22_X1 p10_mult_21_U839 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1388), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1346), .ZN(p10_mult_21_n1328)
         );
  OAI22_X1 p10_mult_21_U840 ( .A1(n904), .A2(p10_mult_21_n1094), .B1(A2[4]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1346) );
  XNOR2_X1 p10_mult_21_U847 ( .A(p10_mult_21_n1392), .B(p10_mult_21_n1385), 
        .ZN(p10_mult_21_n1353) );
  XNOR2_X1 p10_mult_21_U593 ( .A(p10_mult_21_n1105), .B(p10_mult_21_n1103), 
        .ZN(p10_mult_21_n1099) );
  XNOR2_X1 p10_mult_21_U609 ( .A(p10_mult_21_n1101), .B(p10_mult_21_n1102), 
        .ZN(p10_mult_21_n1105) );
  AOI222_X1 p10_mult_21_U616 ( .A1(p10_mult_21_n1134), .A2(p10_mult_21_n1135), 
        .B1(p10_mult_21_n1134), .B2(p10_mult_21_n1136), .C1(p10_mult_21_n1135), 
        .C2(p10_mult_21_n1136), .ZN(p10_mult_21_n1098) );
  AOI222_X1 p10_mult_21_U631 ( .A1(p10_mult_21_n1159), .A2(p10_mult_21_n1160), 
        .B1(p10_mult_21_n1159), .B2(p10_mult_21_n1161), .C1(p10_mult_21_n1160), 
        .C2(p10_mult_21_n1161), .ZN(p10_mult_21_n1136) );
  XNOR2_X1 p10_mult_21_U799 ( .A(p10_mult_21_n1155), .B(p10_mult_21_n1156), 
        .ZN(p10_mult_21_n1367) );
  XNOR2_X1 p10_mult_21_U811 ( .A(p10_mult_21_n1154), .B(p10_mult_21_n1372), 
        .ZN(p10_mult_21_n1160) );
  AOI222_X1 p10_mult_21_U783 ( .A1(p10_mult_21_n1357), .A2(p10_mult_21_n1356), 
        .B1(p10_mult_21_n1357), .B2(p10_mult_21_n1354), .C1(p10_mult_21_n1356), 
        .C2(p10_mult_21_n1354), .ZN(p10_mult_21_n1159) );
  OAI22_X1 p10_mult_21_U784 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1360), 
        .B1(n735), .B2(p10_mult_21_n1361), .ZN(p10_mult_21_n1354) );
  OAI222_X1 p10_mult_21_U786 ( .A1(p10_mult_21_n1343), .A2(p10_mult_21_n1344), 
        .B1(p10_mult_21_n1343), .B2(p10_mult_21_n1342), .C1(p10_mult_21_n1344), 
        .C2(p10_mult_21_n1342), .ZN(p10_mult_21_n1362) );
  OAI22_X1 p10_mult_21_U787 ( .A1(n906), .A2(p10_mult_21_n1363), .B1(
        p10_mult_21_n1294), .B2(p10_mult_21_n1345), .ZN(p10_mult_21_n1342) );
  OAI22_X1 p10_mult_21_U790 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1361), 
        .B1(n735), .B2(p10_mult_21_n1347), .ZN(p10_mult_21_n1344) );
  OAI22_X1 p10_mult_21_U791 ( .A1(p10_mult_21_n1046), .A2(p10_mult_21_n1025), 
        .B1(A2[6]), .B2(reg4[5]), .ZN(p10_mult_21_n1347) );
  OAI22_X1 p10_mult_21_U792 ( .A1(p10_mult_21_n1046), .A2(p10_mult_21_n983), 
        .B1(A2[7]), .B2(reg4[5]), .ZN(p10_mult_21_n1361) );
  OAI22_X1 p10_mult_21_U793 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1364), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1349), .ZN(p10_mult_21_n1343)
         );
  OAI22_X1 p10_mult_21_U794 ( .A1(n901), .A2(p10_mult_21_n1175), .B1(A2[2]), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1349) );
  NOR2_X1 p10_mult_21_U795 ( .A1(p10_mult_21_n1365), .A2(p10_mult_21_n1366), 
        .ZN(p10_mult_21_n1357) );
  AOI21_X1 p10_mult_21_U845 ( .B1(p10_mult_21_n1390), .B2(p10_mult_21_n880), 
        .A(p10_mult_21_n1391), .ZN(p10_mult_21_n1366) );
  XNOR2_X1 p10_mult_21_U632 ( .A(p10_mult_21_n1162), .B(p10_mult_21_n1133), 
        .ZN(p10_mult_21_n1134) );
  XNOR2_X1 p10_mult_21_U638 ( .A(p10_mult_21_n1131), .B(p10_mult_21_n1132), 
        .ZN(p10_mult_21_n1162) );
  AOI222_X1 p10_mult_21_U591 ( .A1(p10_mult_21_n1101), .A2(p10_mult_21_n1102), 
        .B1(p10_mult_21_n1101), .B2(p10_mult_21_n1103), .C1(p10_mult_21_n1102), 
        .C2(p10_mult_21_n1103), .ZN(p10_mult_21_n1033) );
  XNOR2_X1 p10_mult_21_U610 ( .A(p10_mult_21_n1122), .B(p10_mult_21_n1097), 
        .ZN(p10_mult_21_n1102) );
  XNOR2_X1 p10_mult_21_U612 ( .A(p10_mult_21_n1095), .B(p10_mult_21_n1096), 
        .ZN(p10_mult_21_n1122) );
  AOI222_X1 p10_mult_21_U615 ( .A1(p10_mult_21_n1131), .A2(p10_mult_21_n1132), 
        .B1(p10_mult_21_n1131), .B2(p10_mult_21_n1133), .C1(p10_mult_21_n1132), 
        .C2(p10_mult_21_n1133), .ZN(p10_mult_21_n1101) );
  AOI222_X1 p10_mult_21_U639 ( .A1(p10_mult_21_n1168), .A2(p10_mult_21_n1169), 
        .B1(p10_mult_21_n1168), .B2(p10_mult_21_n1170), .C1(p10_mult_21_n1169), 
        .C2(p10_mult_21_n1170), .ZN(p10_mult_21_n1132) );
  XNOR2_X1 p10_mult_21_U824 ( .A(p10_mult_21_n1172), .B(p10_mult_21_n1173), 
        .ZN(p10_mult_21_n1170) );
  AOI222_X1 p10_mult_21_U834 ( .A1(p10_mult_21_n1383), .A2(p10_mult_21_n1384), 
        .B1(p10_mult_21_n1383), .B2(p10_mult_21_n1385), .C1(p10_mult_21_n1384), 
        .C2(p10_mult_21_n1385), .ZN(p10_mult_21_n1169) );
  OAI22_X1 p10_mult_21_U848 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1375), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1388), .ZN(p10_mult_21_n1385)
         );
  AOI22_X1 p10_mult_21_U849 ( .A1(reg4[7]), .A2(p10_mult_21_n1062), .B1(A2[5]), 
        .B2(n904), .ZN(p10_mult_21_n1388) );
  AOI22_X1 p10_mult_21_U866 ( .A1(p10_mult_21_n880), .A2(p10_mult_21_n1371), 
        .B1(p10_mult_21_n881), .B2(p10_mult_21_n1390), .ZN(p10_mult_21_n1386)
         );
  OAI22_X1 p10_mult_21_U867 ( .A1(n902), .A2(A2[1]), .B1(p10_mult_21_n1298), 
        .B2(reg4[11]), .ZN(p10_mult_21_n1390) );
  AOI222_X1 p10_mult_21_U833 ( .A1(p10_mult_21_n1380), .A2(p10_mult_21_n1381), 
        .B1(p10_mult_21_n1380), .B2(p10_mult_21_n1382), .C1(p10_mult_21_n1381), 
        .C2(p10_mult_21_n1382), .ZN(p10_mult_21_n1168) );
  OAI22_X1 p10_mult_21_U876 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1368), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1364), .ZN(p10_mult_21_n1381)
         );
  AOI222_X1 p10_mult_21_U545 ( .A1(p10_mult_21_n1036), .A2(p10_mult_21_n1037), 
        .B1(p10_mult_21_n1036), .B2(p10_mult_21_n1038), .C1(p10_mult_21_n1037), 
        .C2(p10_mult_21_n1038), .ZN(p10_mult_21_n1026) );
  OAI22_X1 p10_mult_21_U577 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1043), 
        .B1(n735), .B2(p10_mult_21_n1083), .ZN(p10_mult_21_n1049) );
  OAI22_X1 p10_mult_21_U580 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n1047), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n1085), .ZN(p10_mult_21_n1048)
         );
  OAI22_X1 p10_mult_21_U583 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1059), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1087), .ZN(p10_mult_21_n1050)
         );
  OAI22_X1 p10_mult_21_U584 ( .A1(n901), .A2(p10_mult_21_n955), .B1(A2[8]), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1059) );
  OAI21_X1 p10_mult_21_U585 ( .B1(p10_mult_21_n1089), .B2(p10_mult_21_n1090), 
        .A(p10_mult_21_n1091), .ZN(p10_mult_21_n1064) );
  OAI22_X1 p10_mult_21_U586 ( .A1(p10_mult_21_n1063), .A2(p10_mult_21_n1061), 
        .B1(p10_mult_21_n1092), .B2(p10_mult_21_n1093), .ZN(p10_mult_21_n1065)
         );
  AOI22_X1 p10_mult_21_U587 ( .A1(reg4[13]), .A2(p10_mult_21_n1094), .B1(A2[4]), .B2(n903), .ZN(p10_mult_21_n1061) );
  AOI222_X1 p10_mult_21_U588 ( .A1(p10_mult_21_n1095), .A2(p10_mult_21_n1096), 
        .B1(p10_mult_21_n1095), .B2(p10_mult_21_n1097), .C1(p10_mult_21_n1096), 
        .C2(p10_mult_21_n1097), .ZN(p10_mult_21_n1054) );
  AOI222_X1 p10_mult_21_U613 ( .A1(p10_mult_21_n1125), .A2(p10_mult_21_n1126), 
        .B1(p10_mult_21_n1125), .B2(p10_mult_21_n1127), .C1(p10_mult_21_n1126), 
        .C2(p10_mult_21_n1127), .ZN(p10_mult_21_n1096) );
  OAI22_X1 p10_mult_21_U633 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1118), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1164), .ZN(p10_mult_21_n1126)
         );
  AOI222_X1 p10_mult_21_U614 ( .A1(p10_mult_21_n1128), .A2(p10_mult_21_n1129), 
        .B1(p10_mult_21_n1128), .B2(p10_mult_21_n1130), .C1(p10_mult_21_n1129), 
        .C2(p10_mult_21_n1130), .ZN(p10_mult_21_n1095) );
  OAI22_X1 p10_mult_21_U643 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1119), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1176), .ZN(p10_mult_21_n1130)
         );
  OAI22_X1 p10_mult_21_U641 ( .A1(p10_mult_21_n1063), .A2(p10_mult_21_n1120), 
        .B1(p10_mult_21_n1092), .B2(p10_mult_21_n1174), .ZN(p10_mult_21_n1129)
         );
  OAI21_X1 p10_mult_21_U825 ( .B1(p10_mult_21_n1174), .B2(p10_mult_21_n1063), 
        .A(p10_mult_21_n1378), .ZN(p10_mult_21_n1173) );
  OAI22_X1 p10_mult_21_U828 ( .A1(n903), .A2(p10_mult_21_n1298), .B1(A2[1]), 
        .B2(reg4[13]), .ZN(p10_mult_21_n1174) );
  AOI221_X1 p10_mult_21_U829 ( .B1(p10_mult_21_n1092), .B2(p10_mult_21_n1063), 
        .C1(p10_mult_21_n1092), .C2(A2[0]), .A(n903), .ZN(p10_mult_21_n1172)
         );
  OAI222_X1 p10_mult_21_U572 ( .A1(p10_mult_21_n1071), .A2(p10_mult_21_n1072), 
        .B1(p10_mult_21_n1071), .B2(p10_mult_21_n1073), .C1(p10_mult_21_n1072), 
        .C2(p10_mult_21_n1073), .ZN(p10_mult_21_n1070) );
  AOI222_X1 p10_mult_21_U573 ( .A1(p10_mult_21_n1074), .A2(p10_mult_21_n1075), 
        .B1(p10_mult_21_n1074), .B2(p10_mult_21_n1066), .C1(p10_mult_21_n1075), 
        .C2(p10_mult_21_n1066), .ZN(p10_mult_21_n1051) );
  OAI22_X1 p10_mult_21_U574 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1042), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1076), .ZN(p10_mult_21_n1053)
         );
  AOI222_X1 p10_mult_21_U576 ( .A1(p10_mult_21_n1077), .A2(p10_mult_21_n1078), 
        .B1(p10_mult_21_n1077), .B2(p10_mult_21_n1079), .C1(p10_mult_21_n1078), 
        .C2(p10_mult_21_n1079), .ZN(p10_mult_21_n1036) );
  OAI22_X1 p10_mult_21_U602 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1087), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1118), .ZN(p10_mult_21_n1073)
         );
  OAI22_X1 p10_mult_21_U634 ( .A1(n901), .A2(p10_mult_21_n1025), .B1(A2[6]), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1118) );
  OAI22_X1 p10_mult_21_U603 ( .A1(n901), .A2(p10_mult_21_n983), .B1(A2[7]), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1087) );
  XNOR2_X1 p10_mult_21_U604 ( .A(p10_mult_21_n1071), .B(p10_mult_21_n1072), 
        .ZN(p10_mult_21_n1117) );
  OAI22_X1 p10_mult_21_U605 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1076), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1119), .ZN(p10_mult_21_n1072)
         );
  OAI22_X1 p10_mult_21_U644 ( .A1(n904), .A2(p10_mult_21_n955), .B1(A2[8]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1119) );
  OAI22_X1 p10_mult_21_U606 ( .A1(n904), .A2(p10_mult_21_n935), .B1(A2[9]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1076) );
  OAI22_X1 p10_mult_21_U607 ( .A1(p10_mult_21_n1063), .A2(p10_mult_21_n1093), 
        .B1(p10_mult_21_n1092), .B2(p10_mult_21_n1120), .ZN(p10_mult_21_n1071)
         );
  OAI22_X1 p10_mult_21_U642 ( .A1(n903), .A2(p10_mult_21_n1175), .B1(A2[2]), 
        .B2(reg4[13]), .ZN(p10_mult_21_n1120) );
  AOI22_X1 p10_mult_21_U595 ( .A1(p10_mult_21_n1021), .A2(p10_mult_21_n1084), 
        .B1(p10_mult_21_n1022), .B2(p10_mult_21_n1111), .ZN(p10_mult_21_n1074)
         );
  AOI22_X1 p10_mult_21_U596 ( .A1(A2[11]), .A2(reg4[5]), .B1(p10_mult_21_n1046), .B2(p10_mult_21_n897), .ZN(p10_mult_21_n1084) );
  OAI21_X1 p10_mult_21_U597 ( .B1(p10_mult_21_n1112), .B2(p10_mult_21_n1113), 
        .A(p10_mult_21_n1114), .ZN(p10_mult_21_n1066) );
  NAND2_X1 p10_mult_21_U598 ( .A1(p10_mult_21_n1089), .A2(p10_mult_21_n1091), 
        .ZN(p10_mult_21_n1114) );
  AOI22_X1 p10_mult_21_U600 ( .A1(p10_mult_21_n880), .A2(p10_mult_21_n1086), 
        .B1(p10_mult_21_n881), .B2(p10_mult_21_n1116), .ZN(p10_mult_21_n1075)
         );
  AOI22_X1 p10_mult_21_U601 ( .A1(reg4[11]), .A2(A2[5]), .B1(p10_mult_21_n1062), .B2(n902), .ZN(p10_mult_21_n1086) );
  AOI222_X1 p10_mult_21_U594 ( .A1(p10_mult_21_n1107), .A2(p10_mult_21_n1108), 
        .B1(p10_mult_21_n1107), .B2(p10_mult_21_n1109), .C1(p10_mult_21_n1108), 
        .C2(p10_mult_21_n1109), .ZN(p10_mult_21_n1077) );
  XNOR2_X1 p10_mult_21_U622 ( .A(p10_mult_21_n1123), .B(p10_mult_21_n1124), 
        .ZN(p10_mult_21_n1109) );
  AOI22_X1 p10_mult_21_U623 ( .A1(p10_mult_21_n880), .A2(p10_mult_21_n1116), 
        .B1(p10_mult_21_n881), .B2(p10_mult_21_n1149), .ZN(p10_mult_21_n1124)
         );
  AOI22_X1 p10_mult_21_U624 ( .A1(reg4[11]), .A2(A2[4]), .B1(p10_mult_21_n1094), .B2(n902), .ZN(p10_mult_21_n1116) );
  AOI22_X1 p10_mult_21_U625 ( .A1(p10_mult_21_n1021), .A2(p10_mult_21_n1111), 
        .B1(p10_mult_21_n1022), .B2(p10_mult_21_n1150), .ZN(p10_mult_21_n1123)
         );
  AOI22_X1 p10_mult_21_U626 ( .A1(A2[10]), .A2(reg4[5]), .B1(p10_mult_21_n1046), .B2(p10_mult_21_n921), .ZN(p10_mult_21_n1111) );
  AOI222_X1 p10_mult_21_U629 ( .A1(p10_mult_21_n1155), .A2(p10_mult_21_n1156), 
        .B1(p10_mult_21_n1155), .B2(p10_mult_21_n1157), .C1(p10_mult_21_n1156), 
        .C2(p10_mult_21_n1157), .ZN(p10_mult_21_n1108) );
  OAI22_X1 p10_mult_21_U797 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1164), 
        .B1(p10_mult_21_n937), .B2(p10_mult_21_n1368), .ZN(p10_mult_21_n1158)
         );
  OAI22_X1 p10_mult_21_U880 ( .A1(n901), .A2(p10_mult_21_n1094), .B1(A2[4]), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1368) );
  AOI22_X1 p10_mult_21_U798 ( .A1(reg4[9]), .A2(p10_mult_21_n1062), .B1(A2[5]), 
        .B2(n901), .ZN(p10_mult_21_n1164) );
  AOI22_X1 p10_mult_21_U800 ( .A1(p10_mult_21_n1021), .A2(p10_mult_21_n1150), 
        .B1(p10_mult_21_n1022), .B2(p10_mult_21_n1369), .ZN(p10_mult_21_n1156)
         );
  OAI22_X1 p10_mult_21_U802 ( .A1(p10_mult_21_n955), .A2(p10_mult_21_n1046), 
        .B1(reg4[5]), .B2(A2[8]), .ZN(p10_mult_21_n1360) );
  OAI22_X1 p10_mult_21_U805 ( .A1(p10_mult_21_n935), .A2(reg4[5]), .B1(
        p10_mult_21_n1046), .B2(A2[9]), .ZN(p10_mult_21_n1150) );
  AOI22_X1 p10_mult_21_U809 ( .A1(p10_mult_21_n880), .A2(p10_mult_21_n1149), 
        .B1(p10_mult_21_n881), .B2(p10_mult_21_n1371), .ZN(p10_mult_21_n1155)
         );
  AOI22_X1 p10_mult_21_U871 ( .A1(reg4[11]), .A2(A2[2]), .B1(p10_mult_21_n1175), .B2(n902), .ZN(p10_mult_21_n1371) );
  OAI222_X1 p10_mult_21_U628 ( .A1(p10_mult_21_n1152), .A2(p10_mult_21_n1153), 
        .B1(p10_mult_21_n1152), .B2(p10_mult_21_n1154), .C1(p10_mult_21_n1153), 
        .C2(p10_mult_21_n1154), .ZN(p10_mult_21_n1151) );
  OAI22_X1 p10_mult_21_U817 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1176), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1375), .ZN(p10_mult_21_n1153)
         );
  OAI22_X1 p10_mult_21_U852 ( .A1(n904), .A2(p10_mult_21_n1025), .B1(A2[6]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1375) );
  AOI22_X1 p10_mult_21_U818 ( .A1(reg4[7]), .A2(p10_mult_21_n983), .B1(A2[7]), 
        .B2(n904), .ZN(p10_mult_21_n1176) );
  OAI22_X1 p10_mult_21_U812 ( .A1(n906), .A2(p10_mult_21_n1373), .B1(
        p10_mult_21_n1294), .B2(p10_mult_21_n1374), .ZN(p10_mult_21_n1152) );
  AOI222_X1 p10_mult_21_U500 ( .A1(p10_mult_21_n970), .A2(p10_mult_21_n971), 
        .B1(p10_mult_21_n970), .B2(p10_mult_21_n972), .C1(p10_mult_21_n971), 
        .C2(p10_mult_21_n972), .ZN(p10_mult_21_n926) );
  XNOR2_X1 p10_mult_21_U505 ( .A(p10_mult_21_n963), .B(p10_mult_21_n981), .ZN(
        p10_mult_21_n972) );
  AOI22_X1 p10_mult_21_U506 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n954), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n982), .ZN(p10_mult_21_n961) );
  OAI22_X1 p10_mult_21_U507 ( .A1(n903), .A2(A2[7]), .B1(p10_mult_21_n983), 
        .B2(reg4[13]), .ZN(p10_mult_21_n954) );
  OAI21_X1 p10_mult_21_U508 ( .B1(p10_mult_21_n984), .B2(p10_mult_21_n985), 
        .A(p10_mult_21_n986), .ZN(p10_mult_21_n946) );
  NAND2_X1 p10_mult_21_U509 ( .A1(p10_mult_21_n951), .A2(p10_mult_21_n953), 
        .ZN(p10_mult_21_n986) );
  AOI22_X1 p10_mult_21_U510 ( .A1(A2[13]), .A2(reg4[7]), .B1(n904), .B2(
        p10_mult_21_n868), .ZN(p10_mult_21_n953) );
  OAI22_X1 p10_mult_21_U511 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n960), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n988), .ZN(p10_mult_21_n963) );
  OAI22_X1 p10_mult_21_U512 ( .A1(n902), .A2(p10_mult_21_n935), .B1(A2[9]), 
        .B2(reg4[11]), .ZN(p10_mult_21_n960) );
  XNOR2_X1 p10_mult_21_U514 ( .A(p10_mult_21_n956), .B(p10_mult_21_n989), .ZN(
        p10_mult_21_n971) );
  XNOR2_X1 p10_mult_21_U515 ( .A(p10_mult_21_n957), .B(p10_mult_21_n958), .ZN(
        p10_mult_21_n989) );
  AOI22_X1 p10_mult_21_U516 ( .A1(p10_mult_21_n917), .A2(p10_mult_21_n966), 
        .B1(p10_mult_21_n918), .B2(p10_mult_21_n990), .ZN(p10_mult_21_n958) );
  OAI22_X1 p10_mult_21_U517 ( .A1(n901), .A2(A2[11]), .B1(p10_mult_21_n897), 
        .B2(reg4[9]), .ZN(p10_mult_21_n966) );
  AOI222_X1 p10_mult_21_U518 ( .A1(p10_mult_21_n991), .A2(p10_mult_21_n992), 
        .B1(p10_mult_21_n991), .B2(p10_mult_21_n993), .C1(p10_mult_21_n992), 
        .C2(p10_mult_21_n993), .ZN(p10_mult_21_n957) );
  AOI222_X1 p10_mult_21_U520 ( .A1(p10_mult_21_n995), .A2(p10_mult_21_n996), 
        .B1(p10_mult_21_n995), .B2(p10_mult_21_n997), .C1(p10_mult_21_n996), 
        .C2(p10_mult_21_n997), .ZN(p10_mult_21_n956) );
  AOI222_X1 p10_mult_21_U522 ( .A1(p10_mult_21_n999), .A2(p10_mult_21_n1000), 
        .B1(p10_mult_21_n999), .B2(p10_mult_21_n1001), .C1(p10_mult_21_n1000), 
        .C2(p10_mult_21_n1001), .ZN(p10_mult_21_n970) );
  OAI21_X1 p10_mult_21_U536 ( .B1(p10_mult_21_n1021), .B2(p10_mult_21_n1022), 
        .A(p10_mult_21_n1023), .ZN(p10_mult_21_n991) );
  XNOR2_X1 p10_mult_21_U537 ( .A(p10_mult_21_n993), .B(p10_mult_21_n994), .ZN(
        p10_mult_21_n1020) );
  AOI22_X1 p10_mult_21_U538 ( .A1(p10_mult_21_n862), .A2(p10_mult_21_n982), 
        .B1(p10_mult_21_n863), .B2(p10_mult_21_n1024), .ZN(p10_mult_21_n994)
         );
  OAI22_X1 p10_mult_21_U567 ( .A1(n903), .A2(A2[5]), .B1(p10_mult_21_n1062), 
        .B2(reg4[13]), .ZN(p10_mult_21_n1024) );
  OAI221_X1 p10_mult_21_U830 ( .B1(n907), .B2(n903), .C1(reg4[12]), .C2(
        reg4[13]), .A(p10_mult_21_n1063), .ZN(p10_mult_21_n1092) );
  AOI22_X1 p10_mult_21_U539 ( .A1(reg4[13]), .A2(A2[6]), .B1(p10_mult_21_n1025), .B2(n903), .ZN(p10_mult_21_n982) );
  OAI22_X1 p10_mult_21_U888 ( .A1(n907), .A2(n902), .B1(reg4[11]), .B2(
        reg4[12]), .ZN(p10_mult_21_n1063) );
  XNOR2_X1 p10_mult_21_U526 ( .A(p10_mult_21_n998), .B(p10_mult_21_n996), .ZN(
        p10_mult_21_n1011) );
  OAI22_X1 p10_mult_21_U527 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n988), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n1012), .ZN(p10_mult_21_n996)
         );
  OAI22_X1 p10_mult_21_U528 ( .A1(n902), .A2(p10_mult_21_n955), .B1(A2[8]), 
        .B2(reg4[11]), .ZN(p10_mult_21_n988) );
  AOI22_X1 p10_mult_21_U529 ( .A1(p10_mult_21_n917), .A2(p10_mult_21_n990), 
        .B1(p10_mult_21_n918), .B2(p10_mult_21_n1013), .ZN(p10_mult_21_n998)
         );
  OAI22_X1 p10_mult_21_U563 ( .A1(n901), .A2(A2[9]), .B1(p10_mult_21_n935), 
        .B2(reg4[9]), .ZN(p10_mult_21_n1013) );
  OAI22_X1 p10_mult_21_U530 ( .A1(n901), .A2(A2[10]), .B1(p10_mult_21_n921), 
        .B2(reg4[9]), .ZN(p10_mult_21_n990) );
  OAI22_X1 p10_mult_21_U531 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n984), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1015), .ZN(p10_mult_21_n997)
         );
  AOI22_X1 p10_mult_21_U532 ( .A1(A2[12]), .A2(n904), .B1(reg4[7]), .B2(
        p10_mult_21_n879), .ZN(p10_mult_21_n984) );
  OAI222_X1 p10_mult_21_U534 ( .A1(p10_mult_21_n1017), .A2(p10_mult_21_n1018), 
        .B1(p10_mult_21_n1017), .B2(p10_mult_21_n1019), .C1(p10_mult_21_n1018), 
        .C2(p10_mult_21_n1019), .ZN(p10_mult_21_n1016) );
  OAI21_X1 p10_mult_21_U551 ( .B1(p10_mult_21_n1043), .B2(n735), .A(
        p10_mult_21_n1045), .ZN(p10_mult_21_n993) );
  NAND2_X1 p10_mult_21_U552 ( .A1(p10_mult_21_n1021), .A2(p10_mult_21_n1023), 
        .ZN(p10_mult_21_n1045) );
  AOI22_X1 p10_mult_21_U553 ( .A1(A2[13]), .A2(reg4[5]), .B1(p10_mult_21_n1046), .B2(p10_mult_21_n868), .ZN(p10_mult_21_n1023) );
  AOI22_X1 p10_mult_21_U579 ( .A1(A2[12]), .A2(p10_mult_21_n1046), .B1(reg4[5]), .B2(p10_mult_21_n879), .ZN(p10_mult_21_n1043) );
  OAI22_X1 p10_mult_21_U554 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n1012), 
        .B1(p10_mult_21_n903), .B2(p10_mult_21_n1047), .ZN(p10_mult_21_n1018)
         );
  OAI22_X1 p10_mult_21_U582 ( .A1(n902), .A2(p10_mult_21_n1025), .B1(A2[6]), 
        .B2(reg4[11]), .ZN(p10_mult_21_n1047) );
  AOI22_X1 p10_mult_21_U555 ( .A1(reg4[11]), .A2(p10_mult_21_n983), .B1(A2[7]), 
        .B2(n902), .ZN(p10_mult_21_n1012) );
  OAI22_X1 p10_mult_21_U549 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1015), 
        .B1(p10_mult_21_n985), .B2(p10_mult_21_n1042), .ZN(p10_mult_21_n1017)
         );
  OAI22_X1 p10_mult_21_U575 ( .A1(n904), .A2(p10_mult_21_n921), .B1(A2[10]), 
        .B2(reg4[7]), .ZN(p10_mult_21_n1042) );
  AOI22_X1 p10_mult_21_U550 ( .A1(A2[11]), .A2(n904), .B1(reg4[7]), .B2(
        p10_mult_21_n897), .ZN(p10_mult_21_n1015) );
  XOR2_X1 p10_mult_21_U984 ( .A(p10_mult_21_n1380), .B(p10_mult_21_n1381), .Z(
        p10_mult_21_n1396) );
  XOR2_X1 p10_mult_21_U983 ( .A(p10_mult_21_n1382), .B(p10_mult_21_n1396), .Z(
        p10_mult_21_n1351) );
  XOR2_X1 p10_mult_21_U982 ( .A(p10_mult_21_n1386), .B(p10_mult_21_n1384), .Z(
        p10_mult_21_n1392) );
  XOR2_X1 p10_mult_21_U981 ( .A(p10_mult_21_n1366), .B(p10_mult_21_n1365), .Z(
        p10_mult_21_n1327) );
  XOR2_X1 p10_mult_21_U980 ( .A(p10_mult_21_n1144), .B(p10_mult_21_n1146), .Z(
        p10_mult_21_n1358) );
  XOR2_X1 p10_mult_21_U979 ( .A(p10_mult_21_n1153), .B(p10_mult_21_n1152), .Z(
        p10_mult_21_n1372) );
  XOR2_X1 p10_mult_21_U978 ( .A(p10_mult_21_n1367), .B(p10_mult_21_n1158), .Z(
        p10_mult_21_n1161) );
  XOR2_X1 p10_mult_21_U977 ( .A(p10_mult_21_n1358), .B(p10_mult_21_n1145), .Z(
        p10_mult_21_n1143) );
  XOR2_X1 p10_mult_21_U976 ( .A(p10_mult_21_n1356), .B(p10_mult_21_n1357), .Z(
        p10_mult_21_n1355) );
  XOR2_X1 p10_mult_21_U975 ( .A(p10_mult_21_n1354), .B(p10_mult_21_n1355), .Z(
        p10_mult_21_n1183) );
  XOR2_X1 p10_mult_21_U974 ( .A(p10_mult_21_n1352), .B(p10_mult_21_n1353), .Z(
        p10_mult_21_n1350) );
  XOR2_X1 p10_mult_21_U973 ( .A(p10_mult_21_n1341), .B(p10_mult_21_n1342), .Z(
        p10_mult_21_n1323) );
  XOR2_X1 p10_mult_21_U972 ( .A(p10_mult_21_n1326), .B(p10_mult_21_n1327), .Z(
        p10_mult_21_n1187) );
  XOR2_X1 p10_mult_21_U971 ( .A(p10_mult_21_n1185), .B(p10_mult_21_n1187), .Z(
        p10_mult_21_n1321) );
  XOR2_X1 p10_mult_21_U970 ( .A(p10_mult_21_n1321), .B(p10_mult_21_n1186), .Z(
        p10_mult_21_n1188) );
  XOR2_X1 p10_mult_21_U969 ( .A(p10_mult_21_n1312), .B(p10_mult_21_n1313), .Z(
        p10_mult_21_n1210) );
  XOR2_X1 p10_mult_21_U968 ( .A(p10_mult_21_n1307), .B(p10_mult_21_n1308), .Z(
        p10_mult_21_n1207) );
  XOR2_X1 p10_mult_21_U967 ( .A(p10_mult_21_n1209), .B(p10_mult_21_n1207), .Z(
        p10_mult_21_n1305) );
  XOR2_X1 p10_mult_21_U965 ( .A(p10_mult_21_n1260), .B(p10_mult_21_n1261), .Z(
        p10_mult_21_n1259) );
  XOR2_X1 p10_mult_21_U963 ( .A(p10_mult_21_n1235), .B(p10_mult_21_n1237), .Z(
        p10_mult_21_n1241) );
  XOR2_X1 p10_mult_21_U962 ( .A(p10_mult_21_n1242), .B(p10_mult_21_n1233), .Z(
        p10_mult_21_n1236) );
  XOR2_X1 p10_mult_21_U961 ( .A(p10_mult_21_n1241), .B(p10_mult_21_n1236), .Z(
        p10_mult_21_n1240) );
  XOR2_X1 p10_mult_21_U960 ( .A(p10_mult_21_n1230), .B(p10_mult_21_n1231), .Z(
        p10_mult_21_n1229) );
  XOR2_X1 p10_mult_21_U957 ( .A(p10_mult_21_n1194), .B(p10_mult_21_n1192), .Z(
        p10_mult_21_n1198) );
  XOR2_X1 p10_mult_21_U956 ( .A(p10_mult_21_n1201), .B(p10_mult_21_n1202), .Z(
        p10_mult_21_n1200) );
  XOR2_X1 p10_mult_21_U955 ( .A(p10_mult_21_n1199), .B(p10_mult_21_n1200), .Z(
        p10_mult_21_n1193) );
  XOR2_X1 p10_mult_21_U954 ( .A(p10_mult_21_n1142), .B(p10_mult_21_n1141), .Z(
        p10_mult_21_n1177) );
  XOR2_X1 p10_mult_21_U953 ( .A(p10_mult_21_n1129), .B(p10_mult_21_n1128), .Z(
        p10_mult_21_n1171) );
  XOR2_X1 p10_mult_21_U952 ( .A(p10_mult_21_n1130), .B(p10_mult_21_n1171), .Z(
        p10_mult_21_n1131) );
  XOR2_X1 p10_mult_21_U951 ( .A(p10_mult_21_n1127), .B(p10_mult_21_n1126), .Z(
        p10_mult_21_n1163) );
  XOR2_X1 p10_mult_21_U950 ( .A(p10_mult_21_n1125), .B(p10_mult_21_n1163), .Z(
        p10_mult_21_n1133) );
  XOR2_X1 p10_mult_21_U949 ( .A(p10_mult_21_n1107), .B(p10_mult_21_n1109), .Z(
        p10_mult_21_n1148) );
  XOR2_X1 p10_mult_21_U948 ( .A(p10_mult_21_n1108), .B(p10_mult_21_n1148), .Z(
        p10_mult_21_n1135) );
  XOR2_X1 p10_mult_21_U947 ( .A(p10_mult_21_n1136), .B(p10_mult_21_n1135), .Z(
        p10_mult_21_n1147) );
  XOR2_X1 p10_mult_21_U946 ( .A(p10_mult_21_n1134), .B(p10_mult_21_n1147), .Z(
        p10_mult_21_n1137) );
  XOR2_X1 p10_mult_21_U945 ( .A(p10_mult_21_n1117), .B(p10_mult_21_n1073), .Z(
        p10_mult_21_n1079) );
  XOR2_X1 p10_mult_21_U944 ( .A(p10_mult_21_n1066), .B(p10_mult_21_n1074), .Z(
        p10_mult_21_n1110) );
  XOR2_X1 p10_mult_21_U943 ( .A(p10_mult_21_n1075), .B(p10_mult_21_n1110), .Z(
        p10_mult_21_n1078) );
  XOR2_X1 p10_mult_21_U942 ( .A(p10_mult_21_n1078), .B(p10_mult_21_n1077), .Z(
        p10_mult_21_n1106) );
  XOR2_X1 p10_mult_21_U941 ( .A(p10_mult_21_n1079), .B(p10_mult_21_n1106), .Z(
        p10_mult_21_n1103) );
  XOR2_X1 p10_mult_21_U940 ( .A(p10_mult_21_n1098), .B(p10_mult_21_n1099), .Z(
        p10_mult_21_n1104) );
  XOR2_X1 p10_mult_21_U939 ( .A(p10_mult_21_n1066), .B(p10_mult_21_n1065), .Z(
        p10_mult_21_n1088) );
  XOR2_X1 p10_mult_21_U938 ( .A(p10_mult_21_n1088), .B(p10_mult_21_n1064), .Z(
        p10_mult_21_n1055) );
  XOR2_X1 p10_mult_21_U937 ( .A(p10_mult_21_n1048), .B(p10_mult_21_n1049), .Z(
        p10_mult_21_n1081) );
  XOR2_X1 p10_mult_21_U936 ( .A(p10_mult_21_n1050), .B(p10_mult_21_n1081), .Z(
        p10_mult_21_n1056) );
  XOR2_X1 p10_mult_21_U935 ( .A(p10_mult_21_n1055), .B(p10_mult_21_n1056), .Z(
        p10_mult_21_n1080) );
  XOR2_X1 p10_mult_21_U934 ( .A(p10_mult_21_n1054), .B(p10_mult_21_n1080), .Z(
        p10_mult_21_n1038) );
  XOR2_X1 p10_mult_21_U933 ( .A(p10_mult_21_n1051), .B(p10_mult_21_n1052), .Z(
        p10_mult_21_n1069) );
  XOR2_X1 p10_mult_21_U932 ( .A(p10_mult_21_n1053), .B(p10_mult_21_n1069), .Z(
        p10_mult_21_n1037) );
  XOR2_X1 p10_mult_21_U931 ( .A(p10_mult_21_n1036), .B(p10_mult_21_n1037), .Z(
        p10_mult_21_n1068) );
  XOR2_X1 p10_mult_21_U930 ( .A(p10_mult_21_n1038), .B(p10_mult_21_n1068), .Z(
        p10_mult_21_n1035) );
  XOR2_X1 p10_mult_21_U929 ( .A(p10_mult_21_n1029), .B(p10_mult_21_n1031), .Z(
        p10_mult_21_n1039) );
  XOR2_X1 p10_mult_21_U927 ( .A(p10_mult_21_n1026), .B(p10_mult_21_n1027), .Z(
        p10_mult_21_n1032) );
  XOR2_X1 p10_mult_21_U926 ( .A(p10_mult_21_n1020), .B(p10_mult_21_n991), .Z(
        p10_mult_21_n1001) );
  XOR2_X1 p10_mult_21_U925 ( .A(p10_mult_21_n997), .B(p10_mult_21_n1011), .Z(
        p10_mult_21_n1000) );
  XOR2_X1 p10_mult_21_U924 ( .A(p10_mult_21_n999), .B(p10_mult_21_n1000), .Z(
        p10_mult_21_n1010) );
  XOR2_X1 p10_mult_21_U923 ( .A(p10_mult_21_n1001), .B(p10_mult_21_n1010), .Z(
        p10_mult_21_n979) );
  XOR2_X1 p10_mult_21_U922 ( .A(p10_mult_21_n977), .B(p10_mult_21_n978), .Z(
        p10_mult_21_n1003) );
  XOR2_X1 p10_mult_21_U921 ( .A(p10_mult_21_n979), .B(p10_mult_21_n1003), .Z(
        p10_mult_21_n976) );
  XOR2_X1 p10_mult_21_U920 ( .A(p10_mult_21_n946), .B(p10_mult_21_n961), .Z(
        p10_mult_21_n981) );
  XOR2_X1 p10_mult_21_U919 ( .A(p10_mult_21_n967), .B(n689), .Z(
        p10_mult_21_n973) );
  XOR2_X1 p10_mult_21_U918 ( .A(p10_mult_21_n941), .B(p10_mult_21_n942), .Z(
        p10_mult_21_n959) );
  XOR2_X1 p10_mult_21_U917 ( .A(p10_mult_21_n943), .B(p10_mult_21_n959), .Z(
        p10_mult_21_n931) );
  XOR2_X1 p10_mult_21_U916 ( .A(p10_mult_21_n950), .B(p10_mult_21_n944), .Z(
        p10_mult_21_n930) );
  XOR2_X1 p10_mult_21_U915 ( .A(p10_mult_21_n929), .B(p10_mult_21_n930), .Z(
        p10_mult_21_n949) );
  XOR2_X1 p10_mult_21_U914 ( .A(p10_mult_21_n931), .B(p10_mult_21_n949), .Z(
        p10_mult_21_n928) );
  XOR2_X1 p10_mult_21_U913 ( .A(p10_mult_21_n900), .B(p10_mult_21_n913), .Z(
        p10_mult_21_n933) );
  XOR2_X1 p10_mult_21_U912 ( .A(p10_mult_21_n907), .B(n697), .Z(
        p10_mult_21_n925) );
  XOR2_X1 p10_mult_21_U911 ( .A(p10_mult_21_n916), .B(p10_mult_21_n898), .Z(
        p10_mult_21_n894) );
  XOR2_X1 p10_mult_21_U910 ( .A(p10_mult_21_n892), .B(p10_mult_21_n893), .Z(
        p10_mult_21_n910) );
  XOR2_X1 p10_mult_21_U909 ( .A(p10_mult_21_n894), .B(p10_mult_21_n910), .Z(
        p10_mult_21_n890) );
  XOR2_X1 p10_mult_21_U908 ( .A(p10_mult_21_n874), .B(p10_mult_21_n886), .Z(
        p10_mult_21_n895) );
  XOR2_X1 p10_mult_21_U907 ( .A(p10_mult_21_n895), .B(p10_mult_21_n887), .Z(
        p10_mult_21_n885) );
  XOR2_X1 p10_mult_21_U906 ( .A(p10_mult_21_n883), .B(n687), .Z(
        p10_mult_21_n888) );
  XOR2_X1 p10_mult_21_U905 ( .A(p10_mult_21_n872), .B(p10_mult_21_n877), .Z(
        p10_mult_21_n871) );
  MUX2_X1 p10_mult_21_U901 ( .A(p10_mult_21_n848), .B(p10_mult_21_n849), .S(
        reg4[0]), .Z(p10_mult_21_n1225) );
  MUX2_X1 p10_mult_21_U899 ( .A(p10_mult_21_n844), .B(p10_mult_21_n845), .S(
        reg4[0]), .Z(p10_mult_21_n1254) );
  MUX2_X1 p10_mult_21_U897 ( .A(p10_mult_21_n840), .B(p10_mult_21_n841), .S(
        reg4[0]), .Z(p10_mult_21_n1278) );
  MUX2_X1 p10_mult_21_U896 ( .A(p10_mult_21_n838), .B(p10_mult_21_n839), .S(
        reg4[0]), .Z(p10_mult_21_n1270) );
  MUX2_X1 p10_mult_21_U895 ( .A(p10_mult_21_n836), .B(p10_mult_21_n837), .S(
        reg4[0]), .Z(p10_mult_21_n1233) );
  OR2_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U1 ( .A1(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_), .A2(reg7[0]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_) );
  XNOR2_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2 ( .A(reg7[0]), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_), .ZN(fb_0_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_1 ( .A(SUB1_N1), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_1_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_), .S(fb_1_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_2 ( .A(SUB1_N2), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_2_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_), .S(fb_2_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_3 ( .A(SUB1_N3), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_3_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_), .S(fb_3_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_4 ( .A(SUB1_N4), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_4_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_), .S(fb_4_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_5 ( .A(SUB1_N5), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_5_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_), .S(fb_5_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_6 ( .A(SUB1_N6), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_6_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_), .S(fb_6_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_7 ( .A(SUB1_N7), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_7_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_), .S(fb_7_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_8 ( .A(SUB1_N8), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_8_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_), .S(fb_8_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_9 ( .A(SUB1_N9), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_9_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_), .S(fb_9_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_10 ( .A(SUB1_N10), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_10_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_), .S(fb_10_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_11 ( .A(SUB1_N11), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_), .S(fb_11_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_12 ( .A(SUB1_N12), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_), .S(fb_12_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_13 ( .A(SUB1_N13), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_13_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_), .S(fb_13_) );
  AND2_X1 s6_add_21_U1 ( .A1(mul1_reg[0]), .A2(mul2_reg[0]), .ZN(
        s6_add_21_carry_1_) );
  XOR2_X1 s6_add_21_U2 ( .A(mul2_reg[0]), .B(mul1_reg[0]), .Z(sig_ff1_0_) );
  FA_X1 s6_add_21_U1_1 ( .A(mul1_reg[1]), .B(mul2_reg[1]), .CI(
        s6_add_21_carry_1_), .CO(s6_add_21_carry_2_), .S(sig_ff1_1_) );
  FA_X1 s6_add_21_U1_2 ( .A(mul1_reg[2]), .B(mul2_reg[2]), .CI(
        s6_add_21_carry_2_), .CO(s6_add_21_carry_3_), .S(sig_ff1_2_) );
  FA_X1 s6_add_21_U1_3 ( .A(mul1_reg[3]), .B(mul2_reg[3]), .CI(
        s6_add_21_carry_3_), .CO(s6_add_21_carry_4_), .S(sig_ff1_3_) );
  FA_X1 s6_add_21_U1_4 ( .A(mul1_reg[4]), .B(mul2_reg[4]), .CI(
        s6_add_21_carry_4_), .CO(s6_add_21_carry_5_), .S(sig_ff1_4_) );
  FA_X1 s6_add_21_U1_5 ( .A(mul1_reg[5]), .B(mul2_reg[5]), .CI(
        s6_add_21_carry_5_), .CO(s6_add_21_carry_6_), .S(sig_ff1_5_) );
  FA_X1 s6_add_21_U1_6 ( .A(mul1_reg[6]), .B(mul2_reg[6]), .CI(
        s6_add_21_carry_6_), .CO(s6_add_21_carry_7_), .S(sig_ff1_6_) );
  FA_X1 s6_add_21_U1_7 ( .A(mul1_reg[7]), .B(mul2_reg[7]), .CI(
        s6_add_21_carry_7_), .CO(s6_add_21_carry_8_), .S(sig_ff1_7_) );
  FA_X1 s6_add_21_U1_8 ( .A(mul1_reg[8]), .B(mul2_reg[8]), .CI(
        s6_add_21_carry_8_), .CO(s6_add_21_carry_9_), .S(sig_ff1_8_) );
  FA_X1 s6_add_21_U1_9 ( .A(mul1_reg[9]), .B(mul2_reg[9]), .CI(
        s6_add_21_carry_9_), .CO(s6_add_21_carry_10_), .S(sig_ff1_9_) );
  FA_X1 s6_add_21_U1_10 ( .A(mul1_reg[10]), .B(mul2_reg[10]), .CI(
        s6_add_21_carry_10_), .CO(s6_add_21_carry_11_), .S(sig_ff1_10_) );
  FA_X1 s6_add_21_U1_11 ( .A(mul1_reg[11]), .B(mul2_reg[11]), .CI(
        s6_add_21_carry_11_), .CO(s6_add_21_carry_12_), .S(sig_ff1_11_) );
  FA_X1 s6_add_21_U1_12 ( .A(mul1_reg[12]), .B(mul2_reg[12]), .CI(
        s6_add_21_carry_12_), .CO(s6_add_21_carry_13_), .S(sig_ff1_12_) );
  FA_X1 s6_add_21_U1_13 ( .A(mul1_reg[13]), .B(mul2_reg[13]), .CI(
        s6_add_21_carry_13_), .S(sig_ff1_13_) );
  AND2_X1 s7_add_21_U1 ( .A1(mul3_reg[0]), .A2(mul4_reg[0]), .ZN(
        s7_add_21_carry_1_) );
  XOR2_X1 s7_add_21_U2 ( .A(mul4_reg[0]), .B(mul3_reg[0]), .Z(sig_ff2_0_) );
  FA_X1 s7_add_21_U1_1 ( .A(mul3_reg[1]), .B(mul4_reg[1]), .CI(
        s7_add_21_carry_1_), .CO(s7_add_21_carry_2_), .S(sig_ff2_1_) );
  FA_X1 s7_add_21_U1_2 ( .A(mul3_reg[2]), .B(mul4_reg[2]), .CI(
        s7_add_21_carry_2_), .CO(s7_add_21_carry_3_), .S(sig_ff2_2_) );
  FA_X1 s7_add_21_U1_3 ( .A(mul3_reg[3]), .B(mul4_reg[3]), .CI(
        s7_add_21_carry_3_), .CO(s7_add_21_carry_4_), .S(sig_ff2_3_) );
  FA_X1 s7_add_21_U1_4 ( .A(mul3_reg[4]), .B(mul4_reg[4]), .CI(
        s7_add_21_carry_4_), .CO(s7_add_21_carry_5_), .S(sig_ff2_4_) );
  FA_X1 s7_add_21_U1_5 ( .A(mul3_reg[5]), .B(mul4_reg[5]), .CI(
        s7_add_21_carry_5_), .CO(s7_add_21_carry_6_), .S(sig_ff2_5_) );
  FA_X1 s7_add_21_U1_6 ( .A(mul3_reg[6]), .B(mul4_reg[6]), .CI(
        s7_add_21_carry_6_), .CO(s7_add_21_carry_7_), .S(sig_ff2_6_) );
  FA_X1 s7_add_21_U1_7 ( .A(mul3_reg[7]), .B(mul4_reg[7]), .CI(
        s7_add_21_carry_7_), .CO(s7_add_21_carry_8_), .S(sig_ff2_7_) );
  FA_X1 s7_add_21_U1_8 ( .A(mul3_reg[8]), .B(mul4_reg[8]), .CI(
        s7_add_21_carry_8_), .CO(s7_add_21_carry_9_), .S(sig_ff2_8_) );
  FA_X1 s7_add_21_U1_9 ( .A(mul3_reg[9]), .B(mul4_reg[9]), .CI(
        s7_add_21_carry_9_), .CO(s7_add_21_carry_10_), .S(sig_ff2_9_) );
  FA_X1 s7_add_21_U1_10 ( .A(mul3_reg[10]), .B(mul4_reg[10]), .CI(
        s7_add_21_carry_10_), .CO(s7_add_21_carry_11_), .S(sig_ff2_10_) );
  FA_X1 s7_add_21_U1_11 ( .A(mul3_reg[11]), .B(mul4_reg[11]), .CI(
        s7_add_21_carry_11_), .CO(s7_add_21_carry_12_), .S(sig_ff2_11_) );
  FA_X1 s7_add_21_U1_12 ( .A(mul3_reg[12]), .B(mul4_reg[12]), .CI(
        s7_add_21_carry_12_), .CO(s7_add_21_carry_13_), .S(sig_ff2_12_) );
  FA_X1 s7_add_21_U1_13 ( .A(mul3_reg[13]), .B(mul4_reg[13]), .CI(
        s7_add_21_carry_13_), .S(sig_ff2_13_) );
  AND2_X1 s8_add_21_U1 ( .A1(sig_ff1_0_), .A2(sig_ff2_0_), .ZN(
        s8_add_21_carry_1_) );
  XOR2_X1 s8_add_21_U2 ( .A(sig_ff2_0_), .B(sig_ff1_0_), .Z(ff[0]) );
  FA_X1 s8_add_21_U1_1 ( .A(sig_ff1_1_), .B(sig_ff2_1_), .CI(
        s8_add_21_carry_1_), .CO(s8_add_21_carry_2_), .S(ff[1]) );
  FA_X1 s8_add_21_U1_2 ( .A(sig_ff1_2_), .B(sig_ff2_2_), .CI(
        s8_add_21_carry_2_), .CO(s8_add_21_carry_3_), .S(ff[2]) );
  FA_X1 s8_add_21_U1_3 ( .A(sig_ff1_3_), .B(sig_ff2_3_), .CI(
        s8_add_21_carry_3_), .CO(s8_add_21_carry_4_), .S(ff[3]) );
  FA_X1 s8_add_21_U1_4 ( .A(sig_ff1_4_), .B(sig_ff2_4_), .CI(
        s8_add_21_carry_4_), .CO(s8_add_21_carry_5_), .S(ff[4]) );
  FA_X1 s8_add_21_U1_5 ( .A(sig_ff1_5_), .B(sig_ff2_5_), .CI(
        s8_add_21_carry_5_), .CO(s8_add_21_carry_6_), .S(ff[5]) );
  FA_X1 s8_add_21_U1_6 ( .A(sig_ff1_6_), .B(sig_ff2_6_), .CI(
        s8_add_21_carry_6_), .CO(s8_add_21_carry_7_), .S(ff[6]) );
  FA_X1 s8_add_21_U1_7 ( .A(sig_ff1_7_), .B(sig_ff2_7_), .CI(
        s8_add_21_carry_7_), .CO(s8_add_21_carry_8_), .S(ff[7]) );
  FA_X1 s8_add_21_U1_8 ( .A(sig_ff1_8_), .B(sig_ff2_8_), .CI(
        s8_add_21_carry_8_), .CO(s8_add_21_carry_9_), .S(ff[8]) );
  FA_X1 s8_add_21_U1_9 ( .A(sig_ff1_9_), .B(sig_ff2_9_), .CI(
        s8_add_21_carry_9_), .CO(s8_add_21_carry_10_), .S(ff[9]) );
  FA_X1 s8_add_21_U1_10 ( .A(sig_ff1_10_), .B(sig_ff2_10_), .CI(
        s8_add_21_carry_10_), .CO(s8_add_21_carry_11_), .S(ff[10]) );
  FA_X1 s8_add_21_U1_11 ( .A(sig_ff1_11_), .B(sig_ff2_11_), .CI(
        s8_add_21_carry_11_), .CO(s8_add_21_carry_12_), .S(ff[11]) );
  FA_X1 s8_add_21_U1_12 ( .A(sig_ff1_12_), .B(sig_ff2_12_), .CI(
        s8_add_21_carry_12_), .CO(s8_add_21_carry_13_), .S(ff[12]) );
  FA_X1 s8_add_21_U1_13 ( .A(sig_ff1_13_), .B(sig_ff2_13_), .CI(
        s8_add_21_carry_13_), .S(ff[13]) );
  AND2_X1 s9_add_21_U1 ( .A1(fb_0_), .A2(xin[0]), .ZN(s9_add_21_carry_1_) );
  FA_X1 s9_add_21_U1_1 ( .A(fb_1_), .B(xin[1]), .CI(s9_add_21_carry_1_), .CO(
        s9_add_21_carry_2_), .S(w[1]) );
  FA_X1 s9_add_21_U1_2 ( .A(fb_2_), .B(xin[2]), .CI(s9_add_21_carry_2_), .CO(
        s9_add_21_carry_3_), .S(w[2]) );
  FA_X1 s9_add_21_U1_3 ( .A(fb_3_), .B(xin[3]), .CI(s9_add_21_carry_3_), .CO(
        s9_add_21_carry_4_), .S(w[3]) );
  FA_X1 s9_add_21_U1_4 ( .A(fb_4_), .B(xin[4]), .CI(s9_add_21_carry_4_), .CO(
        s9_add_21_carry_5_), .S(w[4]) );
  FA_X1 s9_add_21_U1_5 ( .A(fb_5_), .B(xin[5]), .CI(s9_add_21_carry_5_), .CO(
        s9_add_21_carry_6_), .S(w[5]) );
  FA_X1 s9_add_21_U1_6 ( .A(fb_6_), .B(xin[6]), .CI(s9_add_21_carry_6_), .CO(
        s9_add_21_carry_7_), .S(w[6]) );
  FA_X1 s9_add_21_U1_7 ( .A(fb_7_), .B(xin[7]), .CI(s9_add_21_carry_7_), .CO(
        s9_add_21_carry_8_), .S(w[7]) );
  FA_X1 s9_add_21_U1_8 ( .A(fb_8_), .B(xin[8]), .CI(s9_add_21_carry_8_), .CO(
        s9_add_21_carry_9_), .S(w[8]) );
  FA_X1 s9_add_21_U1_9 ( .A(fb_9_), .B(xin[9]), .CI(s9_add_21_carry_9_), .CO(
        s9_add_21_carry_10_), .S(w[9]) );
  FA_X1 s9_add_21_U1_10 ( .A(fb_10_), .B(xin[10]), .CI(s9_add_21_carry_10_), 
        .CO(s9_add_21_carry_11_), .S(w[10]) );
  FA_X1 s9_add_21_U1_11 ( .A(fb_11_), .B(xin[11]), .CI(s9_add_21_carry_11_), 
        .CO(s9_add_21_carry_12_), .S(w[11]) );
  FA_X1 s9_add_21_U1_12 ( .A(fb_12_), .B(xin[12]), .CI(s9_add_21_carry_12_), 
        .CO(s9_add_21_carry_13_), .S(w[12]) );
  FA_X1 s9_add_21_U1_13 ( .A(fb_13_), .B(xin[13]), .CI(s9_add_21_carry_13_), 
        .S(w[13]) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG186_S8 ( .D(REGISTER4_n254), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[12]), .QN(p9_mult_21_n1379) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG159_S14 ( .D(REGISTER4_n260), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[6]), .QN(p9_mult_21_n1393) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG86_S18 ( .D(REGISTER3_n264), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[2]) );
  DFFR_X1 MY_CLK_r_REG202_S1 ( .D(xin_in[9]), .CK(CLK), .RN(RST_n), .Q(n70) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG198_S6 ( .D(REGISTER4_n253), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[13]), .QN(p9_mult_21_n867) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG135_S14 ( .D(REGISTER4_n257), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[9]), .QN(p9_mult_21_n939) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG180_S10 ( .D(REGISTER4_n255), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[11]), .QN(p9_mult_21_n905) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG108_S18 ( .D(REGISTER3_n265), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[1]), .QN(p8_mult_21_n703) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG151_S14 ( .D(REGISTER4_n259), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[7]), .QN(p9_mult_21_n987) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG129_S16 ( .D(REGISTER4_n263), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[3]), .QN(p9_mult_21_n1115) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG126_S15 ( .D(REGISTER3_n263), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[3]), .QN(p8_mult_21_n819) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG167_S14 ( .D(REGISTER4_n261), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[5]), .QN(p9_mult_21_n1046) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG112_S16 ( .D(REGISTER1_n266), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[0]), .QN(p6_mult_21_n692) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG82_S16 ( .D(REGISTER1_n264), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[2]) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG124_S14 ( .D(REGISTER2_n263), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[3]), .QN(p7_mult_21_n1126) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG104_S16 ( .D(REGISTER1_n265), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[1]), .QN(p6_mult_21_n704) );
  DFFR_X1 REG41_MY_CLK_r_REG185_S7 ( .D(REG41_n254), .CK(CLK), .RN(RST_n), .Q(
        reg5[12]) );
  DFFR_X1 REG41_MY_CLK_r_REG172_S11 ( .D(REG41_n256), .CK(CLK), .RN(RST_n), 
        .Q(reg5[10]) );
  DFFR_X1 REG41_MY_CLK_r_REG166_S13 ( .D(REG41_n261), .CK(CLK), .RN(RST_n), 
        .Q(reg5[5]) );
  DFFR_X1 REG41_MY_CLK_r_REG158_S13 ( .D(REG41_n260), .CK(CLK), .RN(RST_n), 
        .Q(reg5[6]) );
  DFFR_X1 REG41_MY_CLK_r_REG142_S13 ( .D(REG41_n258), .CK(CLK), .RN(RST_n), 
        .Q(reg5[8]) );
  DFFR_X1 REG41_MY_CLK_r_REG120_S15 ( .D(REG41_n262), .CK(CLK), .RN(RST_n), 
        .Q(reg5[4]) );
  DFFR_X1 REG41_MY_CLK_r_REG118_S18 ( .D(REG41_n266), .CK(CLK), .RN(RST_n), 
        .Q(reg5[0]) );
  DFFR_X1 REG41_MY_CLK_r_REG88_S18 ( .D(REG41_n264), .CK(CLK), .RN(RST_n), .Q(
        reg5[2]) );
  DFFR_X1 REG41_MY_CLK_r_REG197_S5 ( .D(REG41_n253), .CK(CLK), .RN(RST_n), .Q(
        reg5[13]) );
  DFFR_X1 REG41_MY_CLK_r_REG110_S18 ( .D(REG41_n265), .CK(CLK), .RN(RST_n), 
        .Q(reg5[1]) );
  DFFR_X1 REG41_MY_CLK_r_REG179_S9 ( .D(REG41_n255), .CK(CLK), .RN(RST_n), .Q(
        reg5[11]) );
  DFFR_X1 REG41_MY_CLK_r_REG150_S13 ( .D(REG41_n259), .CK(CLK), .RN(RST_n), 
        .Q(reg5[7]) );
  DFFR_X1 REG41_MY_CLK_r_REG134_S13 ( .D(REG41_n257), .CK(CLK), .RN(RST_n), 
        .Q(reg5[9]) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG89_S19 ( .D(REGISTER4_n264), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[2]), .QN(p9_mult_21_n1394) );
  DFFR_X1 MY_CLK_r_REG211_S1 ( .D(xin_in[3]), .CK(CLK), .RN(RST_n), .Q(n79) );
  DFFR_X1 MY_CLK_r_REG210_S1 ( .D(xin_in[4]), .CK(CLK), .RN(RST_n), .Q(n78) );
  DFFR_X1 MY_CLK_r_REG209_S1 ( .D(xin_in[5]), .CK(CLK), .RN(RST_n), .Q(n77) );
  DFFR_X1 MY_CLK_r_REG208_S1 ( .D(xin_in[6]), .CK(CLK), .RN(RST_n), .Q(n76) );
  DFFR_X1 MY_CLK_r_REG207_S1 ( .D(xin_in[7]), .CK(CLK), .RN(RST_n), .Q(n75) );
  DFFR_X1 MY_CLK_r_REG206_S1 ( .D(xin_in[8]), .CK(CLK), .RN(RST_n), .Q(n74) );
  DFFR_X1 MY_CLK_r_REG205_S1 ( .D(xin_in[0]), .CK(CLK), .RN(RST_n), .Q(n73) );
  DFFR_X1 MY_CLK_r_REG204_S1 ( .D(xin_in[1]), .CK(CLK), .RN(RST_n), .Q(n72) );
  DFFR_X1 MY_CLK_r_REG203_S1 ( .D(xin_in[2]), .CK(CLK), .RN(RST_n), .Q(n71) );
  DFFR_X1 MY_CLK_r_REG201_S1 ( .D(xin_in[10]), .CK(CLK), .RN(RST_n), .Q(n69)
         );
  DFFR_X1 MY_CLK_r_REG200_S1 ( .D(xin_in[11]), .CK(CLK), .RN(RST_n), .Q(n68)
         );
  DFFR_X1 MY_CLK_r_REG199_S1 ( .D(xin_in[12]), .CK(CLK), .RN(RST_n), .Q(n67)
         );
  DFFR_X1 MY_CLK_r_REG1_S1 ( .D(xin_in[13]), .CK(CLK), .RN(RST_n), .Q(n66) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG119_S19 ( .D(REGISTER4_n266), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[0]), .QN(p9_mult_21_n1244) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG173_S12 ( .D(REGISTER4_n256), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[10]), .QN(p9_mult_21_n1395) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG143_S14 ( .D(REGISTER4_n258), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[8]), .QN(p9_mult_21_n1397) );
  DFFR_X1 REGISTER4_MY_CLK_r_REG121_S16 ( .D(REGISTER4_n262), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[4]), .QN(p9_mult_21_n1370) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG183_S7 ( .D(REGISTER3_n254), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[12]) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG170_S11 ( .D(REGISTER3_n256), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[10]) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG156_S13 ( .D(REGISTER3_n260), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[6]) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG140_S13 ( .D(REGISTER3_n258), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[8]) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG116_S18 ( .D(REGISTER3_n266), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[0]), .QN(p8_mult_21_n691) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG52_S15 ( .D(REGISTER3_n262), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[4]) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG181_S6 ( .D(REGISTER2_n254), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[12]), .QN(p7_mult_21_n1386) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG168_S10 ( .D(REGISTER2_n256), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[10]), .QN(p7_mult_21_n1403) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG154_S12 ( .D(REGISTER2_n260), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[6]), .QN(p7_mult_21_n1400) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG138_S12 ( .D(REGISTER2_n258), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[8]), .QN(p7_mult_21_n1331) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG84_S17 ( .D(REGISTER2_n264), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[2]), .QN(p7_mult_21_n1401) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG35_S14 ( .D(REGISTER2_n262), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[4]), .QN(p7_mult_21_n1378) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG114_S17 ( .D(REGISTER2_n266), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[0]), .QN(p7_mult_21_n1260) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG193_S4 ( .D(REGISTER2_n253), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[13]), .QN(p7_mult_21_n876) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG195_S5 ( .D(REGISTER3_n253), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[13]), .QN(p8_mult_21_n814) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG175_S8 ( .D(REGISTER2_n255), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[11]), .QN(p7_mult_21_n911) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG162_S12 ( .D(REGISTER2_n261), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[5]), .QN(p7_mult_21_n1053) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG146_S12 ( .D(REGISTER2_n259), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[7]), .QN(p7_mult_21_n992) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG130_S12 ( .D(REGISTER2_n257), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[9]), .QN(p7_mult_21_n945) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG177_S9 ( .D(REGISTER3_n255), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[11]), .QN(p8_mult_21_n812) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG164_S13 ( .D(REGISTER3_n261), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[5]), .QN(p8_mult_21_n806) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG148_S13 ( .D(REGISTER3_n259), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[7]), .QN(p8_mult_21_n808) );
  DFFR_X1 REGISTER3_MY_CLK_r_REG132_S13 ( .D(REGISTER3_n257), .CK(CLK), .RN(
        RST_n), .Q(reg3_reg[9]), .QN(p8_mult_21_n810) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG122_S13 ( .D(REGISTER1_n263), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[3]), .QN(p6_mult_21_n820) );
  DFFR_X1 REGISTER2_MY_CLK_r_REG106_S17 ( .D(REGISTER2_n265), .CK(CLK), .RN(
        RST_n), .Q(reg2_reg[1]), .QN(p7_mult_21_n1261) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG32_S13 ( .D(REGISTER1_n262), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[4]) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG160_S11 ( .D(REGISTER1_n261), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[5]), .QN(p6_mult_21_n807) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG152_S11 ( .D(REGISTER1_n260), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[6]) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG144_S11 ( .D(REGISTER1_n259), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[7]), .QN(p6_mult_21_n809) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG136_S11 ( .D(REGISTER1_n258), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[8]) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG29_S11 ( .D(REGISTER1_n257), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[9]), .QN(p6_mult_21_n811) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG26_S9 ( .D(REGISTER1_n256), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[10]) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG23_S7 ( .D(REGISTER1_n255), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[11]), .QN(p6_mult_21_n813) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG20_S5 ( .D(REGISTER1_n254), .CK(CLK), .RN(
        RST_n), .Q(reg1_reg[12]) );
  DFFR_X1 REGISTER1_MY_CLK_r_REG2_S3 ( .D(REGISTER1_n253), .CK(CLK), .RN(RST_n), .Q(reg1_reg[13]), .QN(p6_mult_21_n815) );
  DFFR_X1 REG3_1_MY_CLK_r_REG66_S16 ( .D(REG3_1_n267), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[0]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG16_S4 ( .D(REG1_1_n267), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[0]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG65_S16 ( .D(REG3_1_n266), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[1]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG15_S4 ( .D(REG1_1_n266), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[1]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG90_S20 ( .D(REG4_1_n266), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[0]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG91_S20 ( .D(REG4_1_n265), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[1]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG64_S16 ( .D(REG3_1_n265), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[2]) );
  DFFR_X1 REG61_MY_CLK_r_REG28_S10 ( .D(REG61_n265), .CK(CLK), .RN(RST_n), .Q(
        reg7[2]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG14_S4 ( .D(REG1_1_n265), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[2]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG49_S15 ( .D(REG2_1_n269), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[1]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG50_S15 ( .D(REG2_1_n270), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[0]) );
  DFFR_X1 REG51_MY_CLK_r_REG80_S15 ( .D(REG51_n265), .CK(CLK), .RN(RST_n), .Q(
        reg6[1]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_1_) );
  DFFR_X1 REG51_MY_CLK_r_REG81_S15 ( .D(REG51_n266), .CK(CLK), .RN(RST_n), .Q(
        reg6[0]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_) );
  DFFR_X1 REG4_1_MY_CLK_r_REG103_S20 ( .D(REG4_1_n264), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[2]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG63_S16 ( .D(REG3_1_n264), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[3]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG13_S4 ( .D(REG1_1_n264), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[3]) );
  DFFR_X1 REG51_MY_CLK_r_REG79_S15 ( .D(REG51_n264), .CK(CLK), .RN(RST_n), .Q(
        reg6[2]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_2_) );
  DFFR_X1 REG2_1_MY_CLK_r_REG48_S15 ( .D(REG2_1_n268), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[2]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG47_S15 ( .D(REG2_1_n267), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[3]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG62_S16 ( .D(REG3_1_n263), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[4]) );
  DFFR_X1 REG61_MY_CLK_r_REG25_S8 ( .D(REG61_n263), .CK(CLK), .RN(RST_n), .Q(
        reg7[4]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG12_S4 ( .D(REG1_1_n263), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[4]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG102_S20 ( .D(REG4_1_n263), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[3]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG61_S16 ( .D(REG3_1_n262), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[5]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG11_S4 ( .D(REG1_1_n262), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[5]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG60_S16 ( .D(REG3_1_n261), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[6]) );
  DFFR_X1 REG61_MY_CLK_r_REG22_S6 ( .D(REG61_n261), .CK(CLK), .RN(RST_n), .Q(
        reg7[6]) );
  DFFR_X1 REG51_MY_CLK_r_REG78_S15 ( .D(REG51_n263), .CK(CLK), .RN(RST_n), .Q(
        reg6[3]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_3_) );
  DFFR_X1 REG2_1_MY_CLK_r_REG46_S15 ( .D(REG2_1_n266), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[4]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG10_S4 ( .D(REG1_1_n261), .CK(CLK), .RN(RST_n), 
        .Q(mul1_reg[6]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG101_S20 ( .D(REG4_1_n262), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[4]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG45_S15 ( .D(REG2_1_n265), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[5]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG59_S16 ( .D(REG3_1_n260), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[7]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG9_S4 ( .D(REG1_1_n260), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[7]) );
  DFFR_X1 REG51_MY_CLK_r_REG77_S15 ( .D(REG51_n262), .CK(CLK), .RN(RST_n), .Q(
        reg6[4]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_4_) );
  DFFR_X1 REG4_1_MY_CLK_r_REG100_S20 ( .D(REG4_1_n261), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[5]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG8_S4 ( .D(REG1_1_n259), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[8]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG58_S16 ( .D(REG3_1_n259), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[8]) );
  DFFR_X1 REG51_MY_CLK_r_REG76_S15 ( .D(REG51_n261), .CK(CLK), .RN(RST_n), .Q(
        reg6[5]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_5_) );
  DFFR_X1 REG61_MY_CLK_r_REG190_S4 ( .D(REG61_n259), .CK(CLK), .RN(RST_n), .Q(
        reg7[8]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG44_S15 ( .D(REG2_1_n264), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[6]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG43_S15 ( .D(REG2_1_n263), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[7]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG99_S20 ( .D(REG4_1_n260), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[6]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG57_S16 ( .D(REG3_1_n258), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[9]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG7_S4 ( .D(REG1_1_n258), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[9]) );
  DFFR_X1 REG51_MY_CLK_r_REG75_S15 ( .D(REG51_n260), .CK(CLK), .RN(RST_n), .Q(
        reg6[6]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_6_) );
  DFFR_X1 REG4_1_MY_CLK_r_REG98_S20 ( .D(REG4_1_n259), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[7]) );
  DFFR_X1 REG51_MY_CLK_r_REG74_S15 ( .D(REG51_n259), .CK(CLK), .RN(RST_n), .Q(
        reg6[7]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_7_) );
  DFFR_X1 REG3_1_MY_CLK_r_REG56_S16 ( .D(REG3_1_n257), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[10]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG6_S4 ( .D(REG1_1_n257), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[10]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG42_S15 ( .D(REG2_1_n262), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[8]) );
  DFFR_X1 REG61_MY_CLK_r_REG188_S4 ( .D(REG61_n257), .CK(CLK), .RN(RST_n), .Q(
        reg7[10]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG97_S20 ( .D(REG4_1_n258), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[8]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG96_S20 ( .D(REG4_1_n257), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[9]) );
  DFFR_X1 REG3_1_MY_CLK_r_REG55_S16 ( .D(REG3_1_n256), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[11]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG5_S4 ( .D(REG1_1_n256), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[11]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG41_S15 ( .D(REG2_1_n261), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[9]) );
  DFFR_X1 REG51_MY_CLK_r_REG73_S15 ( .D(REG51_n258), .CK(CLK), .RN(RST_n), .Q(
        reg6[8]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_8_) );
  DFFR_X1 REG51_MY_CLK_r_REG72_S15 ( .D(REG51_n257), .CK(CLK), .RN(RST_n), .Q(
        reg6[9]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_9_) );
  DFFR_X1 REG3_1_MY_CLK_r_REG54_S16 ( .D(REG3_1_n255), .CK(CLK), .RN(RST_n), 
        .Q(mul3_reg[12]) );
  DFFR_X1 REG4_1_MY_CLK_r_REG95_S20 ( .D(REG4_1_n256), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[10]) );
  DFFR_X1 REG1_1_MY_CLK_r_REG4_S4 ( .D(REG1_1_n255), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[12]) );
  DFFR_X1 REG61_MY_CLK_r_REG19_S4 ( .D(REG61_n255), .CK(CLK), .RN(RST_n), .Q(
        reg7[12]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG40_S15 ( .D(REG2_1_n260), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[10]) );
  DFFR_X1 REG51_MY_CLK_r_REG71_S15 ( .D(REG51_n256), .CK(CLK), .RN(RST_n), .Q(
        reg6[10]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_10_) );
  DFFR_X1 REG4_1_MY_CLK_r_REG94_S20 ( .D(REG4_1_n255), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[11]) );
  DFFR_X1 REG2_1_MY_CLK_r_REG38_S15 ( .D(REG2_1_n258), .CK(CLK), .RN(RST_n), 
        .Q(mul2_reg[12]) );
  DFFR_X1 REG51_MY_CLK_r_REG68_S15 ( .D(REG51_n253), .CK(CLK), .RN(RST_n), .Q(
        reg6[13]), .QN(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_13_) );
  DFFR_X1 REG4_1_MY_CLK_r_REG92_S20 ( .D(REG4_1_n253), .CK(CLK), .RN(RST_n), 
        .Q(mul4_reg[13]) );
  DFFR_X2 REG11_MY_CLK_r_REG105_S16 ( .D(REG11_n265), .CK(CLK), .RN(RST_n), 
        .Q(reg2[1]), .QN(n888) );
  DFFR_X2 REGISTER4_MY_CLK_r_REG111_S19 ( .D(REGISTER4_n265), .CK(CLK), .RN(
        RST_n), .Q(reg4_reg[1]), .QN(p9_mult_21_n1245) );
  DFFR_X2 REG31_MY_CLK_r_REG109_S17 ( .D(REG31_n265), .CK(CLK), .RN(RST_n), 
        .Q(reg4[1]), .QN(n905) );
  DFFR_X2 REG31_MY_CLK_r_REG127_S14 ( .D(REG31_n263), .CK(CLK), .RN(RST_n), 
        .Q(reg4[3]), .QN(n889) );
  DFFR_X2 REG31_MY_CLK_r_REG165_S12 ( .D(REG31_n261), .CK(CLK), .RN(RST_n), 
        .Q(reg4[5]), .QN(p10_mult_21_n1046) );
  NOR2_X1 U375 ( .A1(n905), .A2(A2[8]), .ZN(n369) );
  INV_X1 U376 ( .A(n461), .ZN(n370) );
  MUX2_X1 U377 ( .A(n370), .B(n369), .S(n462), .Z(p10_mult_21_n1208) );
  NOR2_X1 U378 ( .A1(n905), .A2(A2[9]), .ZN(n371) );
  INV_X1 U379 ( .A(p10_mult_21_n1345), .ZN(n372) );
  MUX2_X1 U380 ( .A(n372), .B(n371), .S(n502), .Z(p10_mult_21_n1335) );
  NOR2_X1 U381 ( .A1(n905), .A2(A2[11]), .ZN(n373) );
  INV_X1 U382 ( .A(p10_mult_21_n1374), .ZN(n374) );
  MUX2_X1 U383 ( .A(n374), .B(n373), .S(n540), .Z(p10_mult_21_n1382) );
  NOR2_X1 U384 ( .A1(p9_mult_21_n1245), .A2(B3[9]), .ZN(n375) );
  INV_X1 U385 ( .A(p9_mult_21_n1345), .ZN(n376) );
  MUX2_X1 U386 ( .A(n376), .B(n375), .S(n542), .Z(p9_mult_21_n1335) );
  NOR2_X1 U387 ( .A1(p9_mult_21_n1245), .A2(B3[6]), .ZN(n377) );
  INV_X1 U388 ( .A(n399), .ZN(n378) );
  MUX2_X1 U389 ( .A(n378), .B(n377), .S(n400), .Z(p9_mult_21_n1233) );
  NOR2_X1 U390 ( .A1(p9_mult_21_n1245), .A2(B3[8]), .ZN(n379) );
  INV_X1 U391 ( .A(n459), .ZN(n380) );
  MUX2_X1 U392 ( .A(n380), .B(n379), .S(n460), .Z(p9_mult_21_n1208) );
  NOR2_X1 U393 ( .A1(p9_mult_21_n1245), .A2(B3[7]), .ZN(n381) );
  INV_X1 U394 ( .A(n433), .ZN(n382) );
  MUX2_X1 U395 ( .A(n382), .B(n381), .S(n434), .Z(p9_mult_21_n1225) );
  NOR2_X1 U396 ( .A1(p9_mult_21_n1245), .A2(B3[11]), .ZN(n383) );
  INV_X1 U397 ( .A(p9_mult_21_n1374), .ZN(n384) );
  MUX2_X1 U398 ( .A(n384), .B(n383), .S(n505), .Z(p9_mult_21_n1382) );
  NOR2_X1 U399 ( .A1(p7_mult_21_n1261), .A2(B1[6]), .ZN(n385) );
  INV_X1 U400 ( .A(n431), .ZN(n386) );
  MUX2_X1 U401 ( .A(n386), .B(n385), .S(n432), .Z(p7_mult_21_n1300) );
  NOR2_X1 U402 ( .A1(p7_mult_21_n1261), .A2(B1[5]), .ZN(n387) );
  INV_X1 U403 ( .A(n401), .ZN(n388) );
  MUX2_X1 U404 ( .A(n388), .B(n387), .S(n402), .Z(p7_mult_21_n1284) );
  NOR2_X1 U405 ( .A1(p7_mult_21_n1261), .A2(B1[8]), .ZN(n389) );
  INV_X1 U406 ( .A(n503), .ZN(n390) );
  MUX2_X1 U407 ( .A(n390), .B(n389), .S(n504), .Z(p7_mult_21_n1328) );
  NOR2_X1 U408 ( .A1(p7_mult_21_n1261), .A2(B1[7]), .ZN(n391) );
  INV_X1 U409 ( .A(n463), .ZN(n392) );
  MUX2_X1 U410 ( .A(n392), .B(n391), .S(n464), .Z(p7_mult_21_n1292) );
  NOR2_X1 U411 ( .A1(p7_mult_21_n1261), .A2(B1[11]), .ZN(n393) );
  INV_X1 U412 ( .A(p7_mult_21_n1381), .ZN(n394) );
  MUX2_X1 U413 ( .A(n394), .B(n393), .S(n541), .Z(p7_mult_21_n1389) );
  INV_X1 U414 ( .A(p10_mult_21_n1044), .ZN(p10_mult_21_n1022) );
  AOI22_X1 U415 ( .A1(reg2_reg[2]), .A2(reg2_reg[1]), .B1(p7_mult_21_n1261), 
        .B2(p7_mult_21_n1401), .ZN(p7_mult_21_n1095) );
  OAI221_X2 U416 ( .B1(p9_mult_21_n1370), .B2(p9_mult_21_n1046), .C1(
        reg4_reg[4]), .C2(reg4_reg[5]), .A(p9_mult_21_n1082), .ZN(
        p9_mult_21_n1044) );
  OAI211_X1 U417 ( .C1(p10_mult_21_n1287), .C2(p10_mult_21_n1089), .A(
        p10_mult_21_n1292), .B(p10_mult_21_n1293), .ZN(n395) );
  OAI221_X1 U418 ( .B1(p10_mult_21_n1090), .B2(p10_mult_21_n1287), .C1(
        p10_mult_21_n1090), .C2(p10_mult_21_n1089), .A(reg4[3]), .ZN(n396) );
  AOI22_X1 U419 ( .A1(n395), .A2(n396), .B1(p10_mult_21_n1284), .B2(
        p10_mult_21_n1283), .ZN(n397) );
  OAI21_X1 U420 ( .B1(p10_mult_21_n1284), .B2(p10_mult_21_n1283), .A(n397), 
        .ZN(n398) );
  OAI21_X1 U421 ( .B1(n395), .B2(n396), .A(n398), .ZN(p10_mult_21_n1279) );
  AOI22_X1 U422 ( .A1(B3[7]), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(
        p9_mult_21_n983), .ZN(n399) );
  INV_X1 U423 ( .A(reg4_reg[0]), .ZN(n400) );
  AOI22_X1 U424 ( .A1(B1[6]), .A2(p7_mult_21_n1261), .B1(reg2_reg[1]), .B2(
        p7_mult_21_n1032), .ZN(n401) );
  INV_X1 U425 ( .A(reg2_reg[0]), .ZN(n402) );
  OAI22_X1 U426 ( .A1(p6_mult_21_n692), .A2(p6_mult_21_n691), .B1(
        p6_mult_21_n689), .B2(p6_mult_21_n690), .ZN(n403) );
  OAI22_X1 U427 ( .A1(p6_mult_21_n707), .A2(p6_mult_21_n708), .B1(
        p6_mult_21_n706), .B2(p6_mult_21_n705), .ZN(n404) );
  NAND3_X1 U428 ( .A1(p6_mult_21_n722), .A2(reg1_reg[3]), .A3(p6_mult_21_n837), 
        .ZN(n405) );
  OAI21_X1 U429 ( .B1(p6_mult_21_n706), .B2(p6_mult_21_n820), .A(n405), .ZN(
        n406) );
  INV_X1 U430 ( .A(n406), .ZN(n407) );
  XNOR2_X1 U431 ( .A(n403), .B(n404), .ZN(n408) );
  AOI222_X1 U432 ( .A1(n407), .A2(p6_mult_21_n839), .B1(n407), .B2(n408), .C1(
        p6_mult_21_n839), .C2(n408), .ZN(n409) );
  OAI211_X1 U433 ( .C1(p6_mult_21_n314), .C2(n409), .A(n403), .B(n404), .ZN(
        n410) );
  NAND2_X1 U434 ( .A1(p6_mult_21_n314), .A2(n409), .ZN(n411) );
  NAND2_X1 U435 ( .A1(n410), .A2(n411), .ZN(p6_mult_21_n681) );
  AOI221_X1 U436 ( .B1(p6_mult_21_n740), .B2(p6_mult_21_n742), .C1(B0[0]), 
        .C2(p6_mult_21_n742), .A(p6_mult_21_n809), .ZN(n412) );
  XNOR2_X1 U437 ( .A(reg1_reg[7]), .B(B0[0]), .ZN(n413) );
  OAI22_X1 U438 ( .A1(p6_mult_21_n742), .A2(n413), .B1(p6_mult_21_n740), .B2(
        p6_mult_21_n743), .ZN(n414) );
  XOR2_X1 U439 ( .A(n412), .B(n414), .Z(p6_mult_21_n304) );
  AND2_X1 U440 ( .A1(n412), .A2(n414), .ZN(p6_mult_21_n303) );
  AOI221_X1 U441 ( .B1(p8_mult_21_n739), .B2(p8_mult_21_n741), .C1(B2[0]), 
        .C2(p8_mult_21_n741), .A(p8_mult_21_n808), .ZN(n415) );
  XNOR2_X1 U442 ( .A(reg3_reg[7]), .B(B2[0]), .ZN(n416) );
  OAI22_X1 U443 ( .A1(p8_mult_21_n741), .A2(n416), .B1(p8_mult_21_n739), .B2(
        p8_mult_21_n742), .ZN(n417) );
  XOR2_X1 U444 ( .A(n415), .B(n417), .Z(p8_mult_21_n304) );
  AND2_X1 U445 ( .A1(n415), .A2(n417), .ZN(p8_mult_21_n303) );
  OAI22_X1 U446 ( .A1(p11_mult_21_n724), .A2(p11_mult_21_n728), .B1(
        p11_mult_21_n727), .B2(p11_mult_21_n726), .ZN(n418) );
  AOI222_X1 U447 ( .A1(p11_mult_21_n311), .A2(p11_mult_21_n308), .B1(
        p11_mult_21_n311), .B2(n418), .C1(p11_mult_21_n308), .C2(n418), .ZN(
        n419) );
  XOR2_X1 U448 ( .A(p11_mult_21_n404), .B(p11_mult_21_n417), .Z(n420) );
  OAI22_X1 U449 ( .A1(p11_mult_21_n682), .A2(p11_mult_21_n313), .B1(n420), 
        .B2(p11_mult_21_n312), .ZN(n421) );
  AOI21_X1 U450 ( .B1(n420), .B2(p11_mult_21_n312), .A(n421), .ZN(n422) );
  AOI21_X1 U451 ( .B1(p11_mult_21_n313), .B2(p11_mult_21_n682), .A(n422), .ZN(
        n423) );
  AOI222_X1 U452 ( .A1(p11_mult_21_n404), .A2(p11_mult_21_n417), .B1(
        p11_mult_21_n404), .B2(p11_mult_21_n312), .C1(p11_mult_21_n417), .C2(
        p11_mult_21_n312), .ZN(n424) );
  XOR2_X1 U453 ( .A(p11_mult_21_n308), .B(p11_mult_21_n311), .Z(n425) );
  AOI22_X1 U454 ( .A1(n423), .A2(n424), .B1(n425), .B2(n418), .ZN(n426) );
  OAI21_X1 U455 ( .B1(n425), .B2(n418), .A(n426), .ZN(n427) );
  OAI21_X1 U456 ( .B1(n423), .B2(n424), .A(n427), .ZN(n428) );
  NOR2_X1 U457 ( .A1(n428), .A2(p11_mult_21_n300), .ZN(n429) );
  NAND2_X1 U458 ( .A1(n428), .A2(p11_mult_21_n300), .ZN(n430) );
  OAI21_X1 U459 ( .B1(n419), .B2(n429), .A(n430), .ZN(p11_mult_21_n636) );
  AOI22_X1 U460 ( .A1(B1[7]), .A2(p7_mult_21_n1261), .B1(reg2_reg[1]), .B2(
        p7_mult_21_n988), .ZN(n431) );
  INV_X1 U461 ( .A(reg2_reg[0]), .ZN(n432) );
  AOI22_X1 U462 ( .A1(B3[8]), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(
        p9_mult_21_n955), .ZN(n433) );
  INV_X1 U463 ( .A(reg4_reg[0]), .ZN(n434) );
  XOR2_X1 U464 ( .A(p10_mult_21_n1274), .B(p10_mult_21_n1275), .Z(n435) );
  OAI222_X1 U465 ( .A1(p10_mult_21_n1265), .A2(p10_mult_21_n1270), .B1(
        p10_mult_21_n1265), .B2(n435), .C1(p10_mult_21_n1270), .C2(n435), .ZN(
        n436) );
  INV_X1 U466 ( .A(n436), .ZN(p10_mult_21_n1256) );
  OR2_X1 U467 ( .A1(p8_mult_21_n703), .A2(B2[1]), .ZN(n437) );
  OAI22_X1 U468 ( .A1(p8_mult_21_n689), .A2(n437), .B1(p8_mult_21_n691), .B2(
        p8_mult_21_n688), .ZN(n438) );
  OAI21_X1 U469 ( .B1(p8_mult_21_n836), .B2(p8_mult_21_n721), .A(n438), .ZN(
        n439) );
  AOI21_X1 U470 ( .B1(p8_mult_21_n721), .B2(n437), .A(n439), .ZN(n440) );
  NAND3_X1 U471 ( .A1(p8_mult_21_n836), .A2(reg3_reg[3]), .A3(p8_mult_21_n721), 
        .ZN(n441) );
  OAI21_X1 U472 ( .B1(p8_mult_21_n819), .B2(p8_mult_21_n705), .A(n441), .ZN(
        n442) );
  AOI222_X1 U473 ( .A1(p8_mult_21_n316), .A2(n440), .B1(p8_mult_21_n316), .B2(
        n442), .C1(n440), .C2(n442), .ZN(p8_mult_21_n832) );
  OAI22_X1 U474 ( .A1(p6_mult_21_n723), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n726), .B2(p6_mult_21_n725), .ZN(n443) );
  AOI222_X1 U475 ( .A1(p6_mult_21_n311), .A2(p6_mult_21_n308), .B1(
        p6_mult_21_n311), .B2(n443), .C1(p6_mult_21_n308), .C2(n443), .ZN(n444) );
  XOR2_X1 U476 ( .A(p6_mult_21_n404), .B(p6_mult_21_n417), .Z(n445) );
  OAI22_X1 U477 ( .A1(p6_mult_21_n681), .A2(p6_mult_21_n313), .B1(n445), .B2(
        p6_mult_21_n312), .ZN(n446) );
  AOI21_X1 U478 ( .B1(n445), .B2(p6_mult_21_n312), .A(n446), .ZN(n447) );
  AOI21_X1 U479 ( .B1(p6_mult_21_n313), .B2(p6_mult_21_n681), .A(n447), .ZN(
        n448) );
  XOR2_X1 U480 ( .A(p6_mult_21_n308), .B(p6_mult_21_n311), .Z(n449) );
  AOI222_X1 U481 ( .A1(p6_mult_21_n404), .A2(p6_mult_21_n417), .B1(
        p6_mult_21_n404), .B2(p6_mult_21_n312), .C1(p6_mult_21_n417), .C2(
        p6_mult_21_n312), .ZN(n450) );
  AOI22_X1 U482 ( .A1(n448), .A2(n450), .B1(n449), .B2(n443), .ZN(n451) );
  OAI21_X1 U483 ( .B1(n449), .B2(n443), .A(n451), .ZN(n452) );
  OAI21_X1 U484 ( .B1(n448), .B2(n450), .A(n452), .ZN(n453) );
  NOR2_X1 U485 ( .A1(n453), .A2(p6_mult_21_n300), .ZN(n454) );
  NAND2_X1 U486 ( .A1(n453), .A2(p6_mult_21_n300), .ZN(n455) );
  OAI21_X1 U487 ( .B1(n444), .B2(n454), .A(n455), .ZN(p6_mult_21_n636) );
  AOI221_X1 U488 ( .B1(p8_mult_21_n756), .B2(p8_mult_21_n758), .C1(B2[0]), 
        .C2(p8_mult_21_n758), .A(p8_mult_21_n810), .ZN(n456) );
  XNOR2_X1 U489 ( .A(reg3_reg[9]), .B(B2[0]), .ZN(n457) );
  OAI22_X1 U490 ( .A1(p8_mult_21_n758), .A2(n457), .B1(p8_mult_21_n756), .B2(
        p8_mult_21_n759), .ZN(n458) );
  XOR2_X1 U491 ( .A(n456), .B(n458), .Z(p8_mult_21_n292) );
  AND2_X1 U492 ( .A1(n456), .A2(n458), .ZN(p8_mult_21_n291) );
  AOI22_X1 U493 ( .A1(B3[9]), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(
        p9_mult_21_n935), .ZN(n459) );
  INV_X1 U494 ( .A(reg4_reg[0]), .ZN(n460) );
  AOI22_X1 U495 ( .A1(A2[9]), .A2(n905), .B1(reg4[1]), .B2(p10_mult_21_n935), 
        .ZN(n461) );
  INV_X1 U496 ( .A(reg4[0]), .ZN(n462) );
  AOI22_X1 U497 ( .A1(B1[8]), .A2(p7_mult_21_n1261), .B1(reg2_reg[1]), .B2(
        p7_mult_21_n962), .ZN(n463) );
  INV_X1 U498 ( .A(reg2_reg[0]), .ZN(n464) );
  OAI22_X1 U499 ( .A1(p8_mult_21_n722), .A2(p8_mult_21_n726), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n724), .ZN(n465) );
  XNOR2_X1 U500 ( .A(p8_mult_21_n308), .B(p8_mult_21_n311), .ZN(n466) );
  XNOR2_X1 U501 ( .A(n466), .B(n465), .ZN(n467) );
  OAI21_X1 U502 ( .B1(p8_mult_21_n417), .B2(p8_mult_21_n404), .A(
        p8_mult_21_n312), .ZN(n468) );
  OAI21_X1 U503 ( .B1(n469), .B2(n470), .A(n468), .ZN(n471) );
  NOR3_X1 U504 ( .A1(p8_mult_21_n643), .A2(p8_mult_21_n644), .A3(
        p8_mult_21_n645), .ZN(n472) );
  XNOR2_X1 U505 ( .A(n470), .B(p8_mult_21_n404), .ZN(n473) );
  XNOR2_X1 U506 ( .A(p8_mult_21_n312), .B(n473), .ZN(n474) );
  INV_X1 U507 ( .A(p8_mult_21_n313), .ZN(n475) );
  AOI222_X1 U508 ( .A1(n472), .A2(n474), .B1(n472), .B2(n475), .C1(n474), .C2(
        n475), .ZN(n476) );
  AOI222_X1 U509 ( .A1(n467), .A2(n471), .B1(n467), .B2(n476), .C1(n471), .C2(
        n476), .ZN(n477) );
  AOI222_X1 U510 ( .A1(p8_mult_21_n308), .A2(p8_mult_21_n311), .B1(
        p8_mult_21_n308), .B2(n465), .C1(p8_mult_21_n311), .C2(n465), .ZN(n478) );
  INV_X1 U511 ( .A(p8_mult_21_n300), .ZN(n479) );
  AOI222_X1 U512 ( .A1(n477), .A2(n478), .B1(n477), .B2(n479), .C1(n478), .C2(
        n479), .ZN(p8_mult_21_n636) );
  INV_X1 U513 ( .A(p8_mult_21_n404), .ZN(n469) );
  INV_X1 U514 ( .A(p8_mult_21_n417), .ZN(n470) );
  AOI221_X1 U515 ( .B1(p8_mult_21_n773), .B2(p8_mult_21_n775), .C1(B2[0]), 
        .C2(p8_mult_21_n775), .A(p8_mult_21_n812), .ZN(n480) );
  XNOR2_X1 U516 ( .A(reg3_reg[11]), .B(B2[0]), .ZN(n481) );
  OAI22_X1 U517 ( .A1(p8_mult_21_n775), .A2(n481), .B1(p8_mult_21_n773), .B2(
        p8_mult_21_n776), .ZN(n482) );
  XOR2_X1 U518 ( .A(n480), .B(n482), .Z(p8_mult_21_n276) );
  AND2_X1 U519 ( .A1(n480), .A2(n482), .ZN(p8_mult_21_n275) );
  AOI221_X1 U520 ( .B1(p11_mult_21_n775), .B2(p11_mult_21_n777), .C1(A1[0]), 
        .C2(p11_mult_21_n777), .A(n883), .ZN(n483) );
  XNOR2_X1 U521 ( .A(reg2[11]), .B(A1[0]), .ZN(n484) );
  OAI22_X1 U522 ( .A1(p11_mult_21_n777), .A2(n484), .B1(p11_mult_21_n775), 
        .B2(p11_mult_21_n778), .ZN(n485) );
  XOR2_X1 U523 ( .A(n483), .B(n485), .Z(p11_mult_21_n276) );
  AND2_X1 U524 ( .A1(n483), .A2(n485), .ZN(p11_mult_21_n275) );
  AOI22_X1 U525 ( .A1(p9_mult_21_n987), .A2(n769), .B1(reg4_reg[7]), .B2(B3[0]), .ZN(n486) );
  INV_X1 U526 ( .A(p9_mult_21_n985), .ZN(n487) );
  INV_X1 U527 ( .A(p9_mult_21_n1318), .ZN(n488) );
  AOI22_X1 U528 ( .A1(n486), .A2(n487), .B1(p9_mult_21_n951), .B2(n488), .ZN(
        p9_mult_21_n1250) );
  AOI22_X1 U529 ( .A1(A2[0]), .A2(reg4[7]), .B1(n904), .B2(p10_mult_21_n1287), 
        .ZN(n489) );
  INV_X1 U530 ( .A(p10_mult_21_n985), .ZN(n490) );
  INV_X1 U531 ( .A(p10_mult_21_n1318), .ZN(n491) );
  AOI22_X1 U532 ( .A1(n489), .A2(n490), .B1(p10_mult_21_n951), .B2(n491), .ZN(
        p10_mult_21_n1250) );
  OAI22_X1 U533 ( .A1(p11_mult_21_n708), .A2(p11_mult_21_n709), .B1(
        p11_mult_21_n706), .B2(p11_mult_21_n707), .ZN(n492) );
  OAI22_X1 U534 ( .A1(p11_mult_21_n693), .A2(p11_mult_21_n692), .B1(
        p11_mult_21_n690), .B2(p11_mult_21_n691), .ZN(n493) );
  XOR2_X1 U535 ( .A(n492), .B(n493), .Z(n494) );
  NAND3_X1 U536 ( .A1(reg2[3]), .A2(p11_mult_21_n838), .A3(p11_mult_21_n723), 
        .ZN(n495) );
  OAI21_X1 U537 ( .B1(p11_mult_21_n707), .B2(n575), .A(n495), .ZN(n496) );
  INV_X1 U538 ( .A(p11_mult_21_n840), .ZN(n497) );
  AOI222_X1 U539 ( .A1(n494), .A2(n496), .B1(n494), .B2(n497), .C1(n496), .C2(
        n497), .ZN(n498) );
  INV_X1 U540 ( .A(p11_mult_21_n314), .ZN(n499) );
  NAND2_X1 U541 ( .A1(n492), .A2(n493), .ZN(n500) );
  AOI222_X1 U542 ( .A1(n498), .A2(n499), .B1(n498), .B2(n500), .C1(n499), .C2(
        n500), .ZN(p11_mult_21_n682) );
  OAI21_X1 U543 ( .B1(p9_mult_21_n909), .B2(p9_mult_21_n908), .A(
        p9_mult_21_n907), .ZN(n501) );
  INV_X1 U544 ( .A(n501), .ZN(n796) );
  INV_X1 U545 ( .A(reg4[0]), .ZN(n502) );
  AOI22_X1 U546 ( .A1(B1[9]), .A2(p7_mult_21_n1261), .B1(reg2_reg[1]), .B2(
        p7_mult_21_n941), .ZN(n503) );
  INV_X1 U547 ( .A(reg2_reg[0]), .ZN(n504) );
  INV_X1 U548 ( .A(reg4_reg[0]), .ZN(n505) );
  AOI221_X1 U549 ( .B1(p6_mult_21_n757), .B2(p6_mult_21_n759), .C1(B0[0]), 
        .C2(p6_mult_21_n759), .A(p6_mult_21_n811), .ZN(n506) );
  XNOR2_X1 U550 ( .A(reg1_reg[9]), .B(B0[0]), .ZN(n507) );
  OAI22_X1 U551 ( .A1(p6_mult_21_n759), .A2(n507), .B1(p6_mult_21_n757), .B2(
        p6_mult_21_n760), .ZN(n508) );
  XOR2_X1 U552 ( .A(n506), .B(n508), .Z(p6_mult_21_n292) );
  AND2_X1 U553 ( .A1(n506), .A2(n508), .ZN(p6_mult_21_n291) );
  AOI221_X1 U554 ( .B1(p11_mult_21_n758), .B2(p11_mult_21_n760), .C1(A1[0]), 
        .C2(p11_mult_21_n760), .A(n884), .ZN(n509) );
  XNOR2_X1 U555 ( .A(reg2[9]), .B(A1[0]), .ZN(n510) );
  OAI22_X1 U556 ( .A1(p11_mult_21_n760), .A2(n510), .B1(p11_mult_21_n758), 
        .B2(p11_mult_21_n761), .ZN(n511) );
  XOR2_X1 U557 ( .A(n509), .B(n511), .Z(p11_mult_21_n292) );
  AND2_X1 U558 ( .A1(n509), .A2(n511), .ZN(p11_mult_21_n291) );
  AOI222_X1 U559 ( .A1(p8_mult_21_n413), .A2(p8_mult_21_n292), .B1(
        p8_mult_21_n413), .B2(p8_mult_21_n297), .C1(p8_mult_21_n292), .C2(
        p8_mult_21_n297), .ZN(n512) );
  OAI222_X1 U560 ( .A1(n513), .A2(p8_mult_21_n282), .B1(n513), .B2(
        p8_mult_21_n280), .C1(p8_mult_21_n282), .C2(p8_mult_21_n280), .ZN(n514) );
  XNOR2_X1 U561 ( .A(p8_mult_21_n413), .B(p8_mult_21_n292), .ZN(n515) );
  XNOR2_X1 U562 ( .A(n515), .B(p8_mult_21_n297), .ZN(n516) );
  XNOR2_X1 U563 ( .A(n516), .B(p8_mult_21_n290), .ZN(n517) );
  XNOR2_X1 U564 ( .A(n517), .B(p8_mult_21_n295), .ZN(n518) );
  OAI21_X1 U565 ( .B1(p8_mult_21_n636), .B2(p8_mult_21_n299), .A(
        p8_mult_21_n294), .ZN(n519) );
  NAND2_X1 U566 ( .A1(n519), .A2(p8_mult_21_n641), .ZN(n520) );
  AOI222_X1 U567 ( .A1(n518), .A2(p8_mult_21_n293), .B1(n518), .B2(n520), .C1(
        p8_mult_21_n293), .C2(n520), .ZN(n521) );
  XNOR2_X1 U568 ( .A(p8_mult_21_n282), .B(n512), .ZN(n522) );
  XNOR2_X1 U569 ( .A(n522), .B(p8_mult_21_n280), .ZN(n523) );
  AOI222_X1 U570 ( .A1(n516), .A2(p8_mult_21_n290), .B1(n516), .B2(
        p8_mult_21_n295), .C1(p8_mult_21_n290), .C2(p8_mult_21_n295), .ZN(n524) );
  AOI222_X1 U571 ( .A1(n521), .A2(n523), .B1(n521), .B2(n524), .C1(n523), .C2(
        n524), .ZN(n525) );
  AOI222_X1 U572 ( .A1(p8_mult_21_n268), .A2(n526), .B1(p8_mult_21_n268), .B2(
        n525), .C1(n526), .C2(n525), .ZN(p8_mult_21_n824) );
  INV_X1 U573 ( .A(n512), .ZN(n513) );
  INV_X1 U574 ( .A(n514), .ZN(n526) );
  NAND4_X1 U575 ( .A1(p10_mult_21_n885), .A2(n685), .A3(n686), .A4(n684), .ZN(
        n527) );
  AND3_X1 U576 ( .A1(p10_mult_21_n871), .A2(n706), .A3(n527), .ZN(n707) );
  OAI21_X1 U577 ( .B1(p7_mult_21_n865), .B2(p7_mult_21_n860), .A(
        p7_mult_21_n864), .ZN(n528) );
  AND2_X1 U578 ( .A1(n528), .A2(n848), .ZN(n846) );
  OAI21_X1 U579 ( .B1(p8_mult_21_n685), .B2(p8_mult_21_n686), .A(
        p8_mult_21_n687), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(p8_mult_21_n162), .ZN(n530) );
  XNOR2_X1 U581 ( .A(p8_mult_21_n136), .B(n530), .ZN(n531) );
  INV_X1 U582 ( .A(VIN), .ZN(n532) );
  AOI22_X1 U583 ( .A1(VIN), .A2(n531), .B1(n915), .B2(n532), .ZN(REG3_1_n254)
         );
  OAI21_X1 U584 ( .B1(p9_mult_21_n1289), .B2(p9_mult_21_n1291), .A(
        p9_mult_21_n1290), .ZN(n533) );
  AND2_X1 U585 ( .A1(n533), .A2(n747), .ZN(p9_mult_21_n1279) );
  AND4_X1 U586 ( .A1(p9_mult_21_n1215), .A2(n742), .A3(n741), .A4(n743), .ZN(
        n744) );
  AOI221_X1 U587 ( .B1(p11_mult_21_n724), .B2(p11_mult_21_n726), .C1(A1[0]), 
        .C2(p11_mult_21_n726), .A(n886), .ZN(n534) );
  XNOR2_X1 U588 ( .A(reg2[5]), .B(A1[0]), .ZN(n535) );
  OAI22_X1 U589 ( .A1(p11_mult_21_n726), .A2(n535), .B1(p11_mult_21_n724), 
        .B2(p11_mult_21_n727), .ZN(n536) );
  XOR2_X1 U590 ( .A(n534), .B(n536), .Z(p11_mult_21_n312) );
  AND2_X1 U591 ( .A1(n534), .A2(n536), .ZN(p11_mult_21_n311) );
  AOI22_X1 U592 ( .A1(n901), .A2(p10_mult_21_n1287), .B1(reg4[9]), .B2(A2[0]), 
        .ZN(n537) );
  INV_X1 U593 ( .A(p10_mult_21_n937), .ZN(n538) );
  INV_X1 U594 ( .A(p10_mult_21_n1340), .ZN(n539) );
  AOI22_X1 U595 ( .A1(n537), .A2(n538), .B1(p10_mult_21_n917), .B2(n539), .ZN(
        p10_mult_21_n1307) );
  AOI222_X1 U596 ( .A1(n682), .A2(p10_mult_21_n1240), .B1(n682), .B2(
        p10_mult_21_n1238), .C1(p10_mult_21_n1240), .C2(p10_mult_21_n1238), 
        .ZN(p10_mult_21_n1220) );
  INV_X1 U597 ( .A(reg4[0]), .ZN(n540) );
  INV_X1 U598 ( .A(reg2_reg[0]), .ZN(n541) );
  INV_X1 U599 ( .A(reg4_reg[0]), .ZN(n542) );
  AOI221_X1 U600 ( .B1(p8_mult_21_n722), .B2(p8_mult_21_n724), .C1(B2[0]), 
        .C2(p8_mult_21_n724), .A(p8_mult_21_n806), .ZN(n543) );
  XNOR2_X1 U601 ( .A(reg3_reg[5]), .B(B2[0]), .ZN(n544) );
  OAI22_X1 U602 ( .A1(p8_mult_21_n724), .A2(n544), .B1(p8_mult_21_n722), .B2(
        p8_mult_21_n725), .ZN(n545) );
  XOR2_X1 U603 ( .A(n543), .B(n545), .Z(p8_mult_21_n312) );
  AND2_X1 U604 ( .A1(n543), .A2(n545), .ZN(p8_mult_21_n311) );
  AOI221_X1 U605 ( .B1(p6_mult_21_n774), .B2(p6_mult_21_n776), .C1(B0[0]), 
        .C2(p6_mult_21_n776), .A(p6_mult_21_n813), .ZN(n546) );
  XNOR2_X1 U606 ( .A(reg1_reg[11]), .B(B0[0]), .ZN(n547) );
  OAI22_X1 U607 ( .A1(p6_mult_21_n776), .A2(n547), .B1(p6_mult_21_n774), .B2(
        p6_mult_21_n777), .ZN(n548) );
  XOR2_X1 U608 ( .A(n546), .B(n548), .Z(p6_mult_21_n276) );
  AND2_X1 U609 ( .A1(n546), .A2(n548), .ZN(p6_mult_21_n275) );
  OAI21_X1 U610 ( .B1(p9_mult_21_n969), .B2(n773), .A(p9_mult_21_n967), .ZN(
        n549) );
  AND2_X1 U611 ( .A1(n549), .A2(n802), .ZN(n768) );
  AND3_X1 U612 ( .A1(p10_mult_21_n976), .A2(n729), .A3(n728), .ZN(n550) );
  AOI221_X1 U613 ( .B1(n695), .B2(p10_mult_21_n974), .C1(p10_mult_21_n976), 
        .C2(p10_mult_21_n974), .A(n550), .ZN(n689) );
  INV_X1 U614 ( .A(p8_mult_21_n657), .ZN(n551) );
  INV_X1 U615 ( .A(p8_mult_21_n246), .ZN(n552) );
  AOI222_X1 U616 ( .A1(p8_mult_21_n824), .A2(p8_mult_21_n825), .B1(
        p8_mult_21_n824), .B2(p8_mult_21_n826), .C1(p8_mult_21_n825), .C2(
        p8_mult_21_n826), .ZN(n553) );
  OAI21_X1 U617 ( .B1(p8_mult_21_n246), .B2(n553), .A(p8_mult_21_n257), .ZN(
        n554) );
  OAI21_X1 U618 ( .B1(n551), .B2(n552), .A(n554), .ZN(p8_mult_21_n148) );
  AOI222_X1 U619 ( .A1(p11_mult_21_n826), .A2(p11_mult_21_n827), .B1(
        p11_mult_21_n826), .B2(p11_mult_21_n828), .C1(p11_mult_21_n827), .C2(
        p11_mult_21_n828), .ZN(n555) );
  OAI21_X1 U620 ( .B1(p11_mult_21_n246), .B2(n555), .A(p11_mult_21_n257), .ZN(
        n556) );
  OAI21_X1 U621 ( .B1(n557), .B2(n558), .A(n556), .ZN(p11_mult_21_n148) );
  INV_X1 U622 ( .A(p11_mult_21_n659), .ZN(n557) );
  INV_X1 U623 ( .A(p11_mult_21_n246), .ZN(n558) );
  AOI222_X1 U624 ( .A1(p10_mult_21_n883), .A2(p10_mult_21_n885), .B1(
        p10_mult_21_n883), .B2(n687), .C1(p10_mult_21_n885), .C2(n688), .ZN(
        n712) );
  NAND2_X1 U625 ( .A1(fb_0_), .A2(xin[0]), .ZN(n559) );
  OAI211_X1 U626 ( .C1(fb_0_), .C2(xin[0]), .A(VIN), .B(n559), .ZN(n288) );
  OAI21_X1 U627 ( .B1(p11_mult_21_n687), .B2(p11_mult_21_n688), .A(
        p11_mult_21_n689), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(p11_mult_21_n162), .ZN(n561) );
  XNOR2_X1 U629 ( .A(p11_mult_21_n136), .B(n561), .ZN(n562) );
  INV_X1 U630 ( .A(VIN), .ZN(n563) );
  AOI22_X1 U631 ( .A1(VIN), .A2(n562), .B1(n914), .B2(n563), .ZN(REG61_n254)
         );
  XOR2_X1 U632 ( .A(p10_mult_21_n861), .B(p10_mult_21_n857), .Z(n564) );
  XNOR2_X1 U633 ( .A(p10_mult_21_n860), .B(n564), .ZN(n565) );
  INV_X1 U634 ( .A(VIN), .ZN(n566) );
  AOI22_X1 U635 ( .A1(VIN), .A2(n565), .B1(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_), .B2(n566), .ZN(
        REG51_n254) );
  AOI222_X1 U636 ( .A1(p7_mult_21_n891), .A2(n828), .B1(p7_mult_21_n891), .B2(
        p7_mult_21_n889), .C1(n828), .C2(p7_mult_21_n889), .ZN(n567) );
  XOR2_X1 U637 ( .A(p7_mult_21_n878), .B(p7_mult_21_n880), .Z(n568) );
  XNOR2_X1 U638 ( .A(n567), .B(n568), .ZN(n569) );
  INV_X1 U639 ( .A(VIN), .ZN(n570) );
  AOI22_X1 U640 ( .A1(VIN), .A2(n569), .B1(n917), .B2(n570), .ZN(REG2_1_n259)
         );
  OAI21_X1 U641 ( .B1(p6_mult_21_n686), .B2(p6_mult_21_n687), .A(
        p6_mult_21_n688), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n571), .B(p6_mult_21_n162), .ZN(n572) );
  XNOR2_X1 U643 ( .A(p6_mult_21_n136), .B(n572), .ZN(n573) );
  INV_X1 U644 ( .A(VIN), .ZN(n574) );
  AOI22_X1 U645 ( .A1(VIN), .A2(n573), .B1(n916), .B2(n574), .ZN(REG1_1_n254)
         );
  INV_X2 U646 ( .A(B3[0]), .ZN(n770) );
  INV_X2 U647 ( .A(B1[0]), .ZN(n830) );
  INV_X2 U648 ( .A(B1[0]), .ZN(n831) );
  INV_X2 U649 ( .A(B3[1]), .ZN(n775) );
  INV_X2 U650 ( .A(B1[4]), .ZN(n841) );
  AND2_X1 U651 ( .A1(n727), .A2(n726), .ZN(p10_mult_21_n1100) );
  AOI222_X2 U652 ( .A1(p7_mult_21_n1183), .A2(p7_mult_21_n1184), .B1(
        p7_mult_21_n1183), .B2(p7_mult_21_n1185), .C1(p7_mult_21_n1184), .C2(
        p7_mult_21_n1185), .ZN(p7_mult_21_n1147) );
  AOI222_X2 U653 ( .A1(p7_mult_21_n1104), .A2(p7_mult_21_n1105), .B1(
        p7_mult_21_n1104), .B2(p7_mult_21_n1106), .C1(p7_mult_21_n1105), .C2(
        p7_mult_21_n1106), .ZN(p7_mult_21_n1040) );
  AOI222_X2 U654 ( .A1(p9_mult_21_n1029), .A2(p9_mult_21_n1030), .B1(
        p9_mult_21_n1029), .B2(p9_mult_21_n1031), .C1(p9_mult_21_n1030), .C2(
        p9_mult_21_n1031), .ZN(p9_mult_21_n974) );
  AOI222_X2 U655 ( .A1(p9_mult_21_n929), .A2(p9_mult_21_n930), .B1(
        p9_mult_21_n929), .B2(p9_mult_21_n931), .C1(p9_mult_21_n930), .C2(
        p9_mult_21_n931), .ZN(p9_mult_21_n907) );
  OAI221_X2 U656 ( .B1(n909), .B2(n904), .C1(reg4[6]), .C2(reg4[7]), .A(
        p10_mult_21_n1014), .ZN(p10_mult_21_n985) );
  AOI221_X1 U657 ( .B1(p7_mult_21_n1028), .B2(B1[0]), .C1(p7_mult_21_n1089), 
        .C2(reg2_reg[4]), .A(p7_mult_21_n1053), .ZN(p7_mult_21_n1277) );
  OAI221_X2 U658 ( .B1(p9_mult_21_n1393), .B2(p9_mult_21_n987), .C1(
        reg4_reg[6]), .C2(reg4_reg[7]), .A(p9_mult_21_n1014), .ZN(
        p9_mult_21_n985) );
  INV_X1 U659 ( .A(p7_mult_21_n943), .ZN(n672) );
  OAI221_X4 U660 ( .B1(p9_mult_21_n1397), .B2(p9_mult_21_n939), .C1(
        reg4_reg[8]), .C2(reg4_reg[9]), .A(p9_mult_21_n964), .ZN(
        p9_mult_21_n937) );
  OAI221_X4 U661 ( .B1(n908), .B2(n901), .C1(reg4[8]), .C2(reg4[9]), .A(
        p10_mult_21_n964), .ZN(p10_mult_21_n937) );
  INV_X1 U662 ( .A(p7_mult_21_n909), .ZN(n673) );
  OAI22_X2 U663 ( .A1(n911), .A2(n905), .B1(reg4[1]), .B2(reg4[2]), .ZN(
        p10_mult_21_n1165) );
  OAI22_X2 U664 ( .A1(n909), .A2(p10_mult_21_n1046), .B1(reg4[5]), .B2(reg4[6]), .ZN(p10_mult_21_n1014) );
  XOR2_X2 U665 ( .A(reg1_reg[12]), .B(p6_mult_21_n813), .Z(p6_mult_21_n791) );
  XOR2_X2 U666 ( .A(reg3_reg[12]), .B(p8_mult_21_n812), .Z(p8_mult_21_n790) );
  XOR2_X2 U667 ( .A(reg2[12]), .B(n883), .Z(p11_mult_21_n792) );
  XNOR2_X2 U668 ( .A(reg2[4]), .B(reg2[3]), .ZN(p11_mult_21_n724) );
  XOR2_X2 U669 ( .A(reg1_reg[10]), .B(p6_mult_21_n811), .Z(p6_mult_21_n774) );
  XOR2_X2 U670 ( .A(reg3_reg[10]), .B(p8_mult_21_n810), .Z(p8_mult_21_n773) );
  XOR2_X2 U671 ( .A(reg2[10]), .B(n884), .Z(p11_mult_21_n775) );
  XOR2_X2 U672 ( .A(reg1_reg[8]), .B(p6_mult_21_n809), .Z(p6_mult_21_n757) );
  XOR2_X2 U673 ( .A(reg1_reg[6]), .B(p6_mult_21_n807), .Z(p6_mult_21_n740) );
  XOR2_X2 U674 ( .A(reg3_reg[8]), .B(p8_mult_21_n808), .Z(p8_mult_21_n756) );
  XOR2_X2 U675 ( .A(reg3_reg[6]), .B(p8_mult_21_n806), .Z(p8_mult_21_n739) );
  XOR2_X2 U676 ( .A(reg2[8]), .B(n885), .Z(p11_mult_21_n758) );
  XOR2_X2 U677 ( .A(reg2[6]), .B(n886), .Z(p11_mult_21_n741) );
  XOR2_X2 U678 ( .A(reg1_reg[4]), .B(p6_mult_21_n820), .Z(p6_mult_21_n723) );
  XOR2_X2 U679 ( .A(reg3_reg[4]), .B(p8_mult_21_n819), .Z(p8_mult_21_n722) );
  AOI22_X1 U680 ( .A1(reg4[1]), .A2(p10_mult_21_n1121), .B1(A2[3]), .B2(n905), 
        .ZN(p10_mult_21_n1296) );
  NAND2_X1 U681 ( .A1(n906), .A2(reg4[1]), .ZN(p10_mult_21_n1294) );
  AOI22_X1 U682 ( .A1(reg4[1]), .A2(p10_mult_21_n1175), .B1(A2[2]), .B2(n905), 
        .ZN(p10_mult_21_n1295) );
  AOI22_X1 U683 ( .A1(reg4[1]), .A2(p10_mult_21_n1094), .B1(A2[4]), .B2(n905), 
        .ZN(p10_mult_21_n1286) );
  OAI21_X1 U684 ( .B1(p10_mult_21_n1288), .B2(p10_mult_21_n1165), .A(
        p10_mult_21_n1297), .ZN(p10_mult_21_n1283) );
  OAI22_X1 U685 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1273), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1288), .ZN(p10_mult_21_n1277) );
  AOI22_X1 U686 ( .A1(A2[6]), .A2(n905), .B1(reg4[1]), .B2(p10_mult_21_n1025), 
        .ZN(p10_mult_21_n1303) );
  AOI22_X1 U687 ( .A1(A2[5]), .A2(n905), .B1(reg4[1]), .B2(p10_mult_21_n1062), 
        .ZN(p10_mult_21_n1271) );
  OAI22_X1 U688 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1249), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1272), .ZN(p10_mult_21_n1253) );
  OAI22_X1 U689 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1272), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1273), .ZN(p10_mult_21_n1265) );
  AOI22_X1 U690 ( .A1(A2[8]), .A2(n905), .B1(reg4[1]), .B2(p10_mult_21_n955), 
        .ZN(p10_mult_21_n1310) );
  AOI22_X1 U691 ( .A1(A2[7]), .A2(n905), .B1(reg4[1]), .B2(p10_mult_21_n983), 
        .ZN(p10_mult_21_n1243) );
  OAI22_X1 U692 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1248), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1249), .ZN(p10_mult_21_n1232) );
  OAI22_X1 U693 ( .A1(p10_mult_21_n921), .A2(n905), .B1(reg4[1]), .B2(A2[10]), 
        .ZN(p10_mult_21_n1345) );
  OAI22_X1 U694 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1316), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1248), .ZN(p10_mult_21_n1228) );
  OAI22_X1 U695 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1331), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1316), .ZN(p10_mult_21_n1313) );
  OAI22_X1 U696 ( .A1(p10_mult_21_n897), .A2(n905), .B1(reg4[1]), .B2(A2[11]), 
        .ZN(p10_mult_21_n1363) );
  OAI22_X1 U697 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1348), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1331), .ZN(p10_mult_21_n1206) );
  OAI22_X1 U698 ( .A1(p10_mult_21_n879), .A2(n905), .B1(reg4[1]), .B2(A2[12]), 
        .ZN(p10_mult_21_n1374) );
  OAI22_X1 U699 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1376), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1389), .ZN(p10_mult_21_n1384) );
  AOI22_X1 U700 ( .A1(A2[13]), .A2(reg4[1]), .B1(n905), .B2(p10_mult_21_n868), 
        .ZN(p10_mult_21_n1167) );
  OAI22_X1 U701 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1389), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1348), .ZN(p10_mult_21_n1329) );
  OAI22_X1 U702 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1166), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1376), .ZN(p10_mult_21_n1154) );
  OAI22_X1 U703 ( .A1(p10_mult_21_n1165), .A2(p10_mult_21_n1112), .B1(
        p10_mult_21_n1113), .B2(p10_mult_21_n1166), .ZN(p10_mult_21_n1127) );
  OAI21_X1 U704 ( .B1(reg4[1]), .B2(reg4[0]), .A(p10_mult_21_n1167), .ZN(
        p10_mult_21_n1125) );
  XNOR2_X1 U705 ( .A(p10_mult_21_n1033), .B(p10_mult_21_n1034), .ZN(
        p10_mult_21_n1067) );
  XNOR2_X1 U706 ( .A(p10_mult_21_n906), .B(n681), .ZN(temp5[9]) );
  XNOR2_X1 U707 ( .A(p10_mult_21_n1140), .B(p10_mult_21_n1138), .ZN(temp5[1])
         );
  AOI222_X1 U708 ( .A1(p10_mult_21_n1213), .A2(p10_mult_21_n1214), .B1(
        p10_mult_21_n1213), .B2(p10_mult_21_n1215), .C1(p10_mult_21_n1214), 
        .C2(p10_mult_21_n1215), .ZN(p10_mult_21_n1195) );
  OAI22_X1 U709 ( .A1(n889), .A2(p10_mult_21_n1175), .B1(A2[2]), .B2(reg4[3]), 
        .ZN(p10_mult_21_n1273) );
  AOI222_X1 U710 ( .A1(p10_mult_21_n1220), .A2(p10_mult_21_n1221), .B1(
        p10_mult_21_n1220), .B2(p10_mult_21_n1222), .C1(p10_mult_21_n1222), 
        .C2(p10_mult_21_n1221), .ZN(p10_mult_21_n1214) );
  AOI222_X1 U711 ( .A1(p10_mult_21_n1188), .A2(p10_mult_21_n1189), .B1(
        p10_mult_21_n1188), .B2(p10_mult_21_n1190), .C1(p10_mult_21_n1189), 
        .C2(p10_mult_21_n1190), .ZN(p10_mult_21_n1178) );
  AOI222_X1 U712 ( .A1(p10_mult_21_n1195), .A2(p10_mult_21_n1196), .B1(
        p10_mult_21_n1195), .B2(p10_mult_21_n1197), .C1(p10_mult_21_n1196), 
        .C2(p10_mult_21_n1197), .ZN(p10_mult_21_n1189) );
  XNOR2_X1 U713 ( .A(p10_mult_21_n1250), .B(p10_mult_21_n1251), .ZN(
        p10_mult_21_n1237) );
  NOR2_X1 U714 ( .A1(A2[2]), .A2(n905), .ZN(p10_mult_21_n842) );
  OAI21_X1 U715 ( .B1(A2[1]), .B2(n905), .A(p10_mult_21_n1287), .ZN(
        p10_mult_21_n1292) );
  NOR2_X1 U716 ( .A1(A2[3]), .A2(n905), .ZN(p10_mult_21_n840) );
  NOR2_X1 U717 ( .A1(A2[5]), .A2(n905), .ZN(p10_mult_21_n844) );
  NOR2_X1 U718 ( .A1(A2[4]), .A2(n905), .ZN(p10_mult_21_n838) );
  NOR2_X1 U719 ( .A1(A2[7]), .A2(n905), .ZN(p10_mult_21_n848) );
  NOR2_X1 U720 ( .A1(A2[6]), .A2(n905), .ZN(p10_mult_21_n836) );
  XNOR2_X1 U721 ( .A(n696), .B(p10_mult_21_n974), .ZN(p10_mult_21_n1002) );
  XOR2_X1 U722 ( .A(p10_mult_21_n1219), .B(p10_mult_21_n1216), .Z(n674) );
  XNOR2_X1 U723 ( .A(n674), .B(p10_mult_21_n1217), .ZN(p10_mult_21_n1222) );
  AOI222_X1 U724 ( .A1(p10_mult_21_n1276), .A2(p10_mult_21_n1277), .B1(
        p10_mult_21_n1276), .B2(p10_mult_21_n1278), .C1(p10_mult_21_n1277), 
        .C2(p10_mult_21_n1278), .ZN(p10_mult_21_n1267) );
  AOI222_X1 U725 ( .A1(p10_mult_21_n1258), .A2(p10_mult_21_n1261), .B1(
        p10_mult_21_n1258), .B2(p10_mult_21_n1260), .C1(p10_mult_21_n1261), 
        .C2(p10_mult_21_n1260), .ZN(p10_mult_21_n1238) );
  NOR3_X1 U726 ( .A1(n680), .A2(n679), .A3(n678), .ZN(p10_mult_21_n1255) );
  AOI22_X1 U727 ( .A1(p10_mult_21_n1279), .A2(p10_mult_21_n1280), .B1(
        p10_mult_21_n1283), .B2(p10_mult_21_n1284), .ZN(p10_mult_21_n1282) );
  NOR2_X1 U728 ( .A1(p10_mult_21_n1275), .A2(n694), .ZN(p10_mult_21_n1261) );
  OAI221_X1 U729 ( .B1(p10_mult_21_n1022), .B2(p10_mult_21_n1021), .C1(
        p10_mult_21_n1022), .C2(p10_mult_21_n1287), .A(reg4[5]), .ZN(
        p10_mult_21_n1275) );
  AOI222_X1 U730 ( .A1(p10_mult_21_n907), .A2(n697), .B1(p10_mult_21_n907), 
        .B2(p10_mult_21_n909), .C1(n697), .C2(p10_mult_21_n909), .ZN(n681) );
  NOR3_X1 U731 ( .A1(n677), .A2(n676), .A3(n675), .ZN(n682) );
  AOI22_X1 U732 ( .A1(reg4[3]), .A2(p10_mult_21_n1298), .B1(A2[1]), .B2(n889), 
        .ZN(p10_mult_21_n1288) );
  AOI22_X1 U733 ( .A1(reg4[3]), .A2(p10_mult_21_n1062), .B1(A2[5]), .B2(n889), 
        .ZN(p10_mult_21_n1248) );
  OAI22_X1 U734 ( .A1(p10_mult_21_n1025), .A2(n889), .B1(reg4[3]), .B2(A2[6]), 
        .ZN(p10_mult_21_n1316) );
  OAI22_X1 U735 ( .A1(p10_mult_21_n983), .A2(n889), .B1(reg4[3]), .B2(A2[7]), 
        .ZN(p10_mult_21_n1331) );
  OAI22_X1 U736 ( .A1(p10_mult_21_n955), .A2(n889), .B1(reg4[3]), .B2(A2[8]), 
        .ZN(p10_mult_21_n1348) );
  AOI22_X1 U737 ( .A1(A2[9]), .A2(n889), .B1(reg4[3]), .B2(p10_mult_21_n935), 
        .ZN(p10_mult_21_n1389) );
  OAI22_X1 U738 ( .A1(p10_mult_21_n921), .A2(n889), .B1(reg4[3]), .B2(A2[10]), 
        .ZN(p10_mult_21_n1376) );
  AOI22_X1 U739 ( .A1(A2[11]), .A2(n889), .B1(reg4[3]), .B2(p10_mult_21_n897), 
        .ZN(p10_mult_21_n1166) );
  AOI22_X1 U740 ( .A1(A2[13]), .A2(reg4[3]), .B1(n889), .B2(p10_mult_21_n868), 
        .ZN(p10_mult_21_n1091) );
  AOI22_X1 U741 ( .A1(A2[12]), .A2(n889), .B1(reg4[3]), .B2(p10_mult_21_n879), 
        .ZN(p10_mult_21_n1112) );
  OAI22_X1 U742 ( .A1(n889), .A2(p10_mult_21_n1094), .B1(A2[4]), .B2(reg4[3]), 
        .ZN(p10_mult_21_n1249) );
  OAI22_X1 U743 ( .A1(n889), .A2(p10_mult_21_n1121), .B1(A2[3]), .B2(reg4[3]), 
        .ZN(p10_mult_21_n1272) );
  OAI221_X1 U744 ( .B1(reg4[3]), .B2(A2[0]), .C1(n889), .C2(p10_mult_21_n1287), 
        .A(p10_mult_21_n1090), .ZN(p10_mult_21_n1297) );
  NOR2_X1 U745 ( .A1(p10_mult_21_n1082), .A2(p10_mult_21_n1287), .ZN(
        p10_mult_21_n1276) );
  NOR2_X1 U746 ( .A1(p10_mult_21_n1014), .A2(p10_mult_21_n1287), .ZN(
        p10_mult_21_n1252) );
  OAI221_X1 U747 ( .B1(p10_mult_21_n952), .B2(p10_mult_21_n951), .C1(
        p10_mult_21_n952), .C2(p10_mult_21_n1287), .A(reg4[7]), .ZN(
        p10_mult_21_n1251) );
  NOR2_X1 U748 ( .A1(p10_mult_21_n911), .A2(p10_mult_21_n1287), .ZN(
        p10_mult_21_n1337) );
  NOR2_X1 U749 ( .A1(p10_mult_21_n964), .A2(p10_mult_21_n1287), .ZN(
        p10_mult_21_n1227) );
  OAI221_X1 U750 ( .B1(p10_mult_21_n918), .B2(p10_mult_21_n917), .C1(
        p10_mult_21_n918), .C2(p10_mult_21_n1287), .A(reg4[9]), .ZN(
        p10_mult_21_n1308) );
  OAI221_X1 U751 ( .B1(p10_mult_21_n881), .B2(p10_mult_21_n880), .C1(
        p10_mult_21_n881), .C2(p10_mult_21_n1287), .A(reg4[11]), .ZN(
        p10_mult_21_n1365) );
  NOR2_X1 U752 ( .A1(p10_mult_21_n1063), .A2(p10_mult_21_n1287), .ZN(
        p10_mult_21_n1380) );
  AOI22_X1 U753 ( .A1(reg4[5]), .A2(p10_mult_21_n1121), .B1(A2[3]), .B2(
        p10_mult_21_n1046), .ZN(p10_mult_21_n1246) );
  XNOR2_X1 U754 ( .A(p10_mult_21_n1274), .B(p10_mult_21_n1275), .ZN(
        p10_mult_21_n1264) );
  XNOR2_X1 U755 ( .A(p10_mult_21_n1264), .B(p10_mult_21_n1265), .ZN(
        p10_mult_21_n1269) );
  NAND2_X1 U756 ( .A1(p10_mult_21_n889), .A2(p10_mult_21_n890), .ZN(n686) );
  XNOR2_X1 U757 ( .A(p10_mult_21_n1285), .B(p10_mult_21_n1278), .ZN(
        p10_mult_21_n1280) );
  NAND2_X1 U758 ( .A1(n690), .A2(p10_mult_21_n1281), .ZN(p10_mult_21_n1266) );
  XNOR2_X1 U759 ( .A(p10_mult_21_n926), .B(p10_mult_21_n927), .ZN(
        p10_mult_21_n948) );
  XNOR2_X1 U760 ( .A(p10_mult_21_n980), .B(p10_mult_21_n972), .ZN(
        p10_mult_21_n969) );
  AOI22_X1 U761 ( .A1(reg4[13]), .A2(p10_mult_21_n1121), .B1(A2[3]), .B2(n903), 
        .ZN(p10_mult_21_n1093) );
  OAI22_X1 U762 ( .A1(n902), .A2(A2[3]), .B1(p10_mult_21_n1121), .B2(reg4[11]), 
        .ZN(p10_mult_21_n1149) );
  AOI22_X1 U763 ( .A1(reg4[9]), .A2(p10_mult_21_n1121), .B1(A2[3]), .B2(n901), 
        .ZN(p10_mult_21_n1364) );
  OAI22_X1 U764 ( .A1(n904), .A2(p10_mult_21_n1121), .B1(A2[3]), .B2(reg4[7]), 
        .ZN(p10_mult_21_n1333) );
  NAND2_X1 U765 ( .A1(n691), .A2(n692), .ZN(p10_mult_21_n1284) );
  NAND2_X1 U766 ( .A1(p10_mult_21_n843), .A2(reg4[0]), .ZN(n691) );
  NAND2_X1 U767 ( .A1(p10_mult_21_n842), .A2(n906), .ZN(n692) );
  XNOR2_X1 U768 ( .A(p10_mult_21_n1269), .B(p10_mult_21_n1270), .ZN(
        p10_mult_21_n1268) );
  AOI22_X1 U769 ( .A1(reg4[5]), .A2(A2[1]), .B1(p10_mult_21_n1298), .B2(
        p10_mult_21_n1046), .ZN(p10_mult_21_n1300) );
  NOR2_X1 U770 ( .A1(n693), .A2(p10_mult_21_n1301), .ZN(p10_mult_21_n1274) );
  NOR2_X1 U771 ( .A1(n693), .A2(p10_mult_21_n1301), .ZN(n694) );
  AOI222_X1 U772 ( .A1(p10_mult_21_n1026), .A2(p10_mult_21_n1027), .B1(
        p10_mult_21_n1026), .B2(p10_mult_21_n1028), .C1(p10_mult_21_n1027), 
        .C2(p10_mult_21_n1028), .ZN(n695) );
  XNOR2_X1 U773 ( .A(p10_mult_21_n1277), .B(p10_mult_21_n1276), .ZN(
        p10_mult_21_n1285) );
  XNOR2_X1 U774 ( .A(p10_mult_21_n1100), .B(p10_mult_21_n1104), .ZN(temp5[2])
         );
  XNOR2_X1 U775 ( .A(n704), .B(n703), .ZN(temp5[13]) );
  OAI21_X1 U776 ( .B1(p10_mult_21_n861), .B2(p10_mult_21_n860), .A(n700), .ZN(
        n699) );
  OAI21_X1 U777 ( .B1(n701), .B2(n700), .A(n699), .ZN(n704) );
  NAND2_X1 U778 ( .A1(n687), .A2(p10_mult_21_n885), .ZN(n705) );
  NAND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n688), .A2(p10_mult_21_n883), .ZN(n708) );
  NAND3_X1 U781 ( .A1(n708), .A2(n705), .A3(n734), .ZN(n711) );
  FA_X1 U782 ( .A(p10_mult_21_n871), .B(p10_mult_21_n869), .CI(n712), .S(
        temp5[11]) );
  NAND2_X1 U783 ( .A1(p10_mult_21_n908), .A2(p10_mult_21_n909), .ZN(n718) );
  OAI21_X1 U784 ( .B1(p10_mult_21_n908), .B2(p10_mult_21_n909), .A(
        p10_mult_21_n907), .ZN(n719) );
  NAND3_X1 U785 ( .A1(n719), .A2(p10_mult_21_n890), .A3(n718), .ZN(n684) );
  AOI222_X1 U786 ( .A1(p10_mult_21_n926), .A2(p10_mult_21_n927), .B1(
        p10_mult_21_n926), .B2(p10_mult_21_n928), .C1(p10_mult_21_n927), .C2(
        p10_mult_21_n928), .ZN(n683) );
  NAND2_X1 U787 ( .A1(n689), .A2(p10_mult_21_n967), .ZN(n722) );
  NAND2_X1 U788 ( .A1(p10_mult_21_n968), .A2(p10_mult_21_n969), .ZN(n720) );
  NAND2_X1 U789 ( .A1(p10_mult_21_n967), .A2(p10_mult_21_n969), .ZN(n721) );
  AOI222_X1 U790 ( .A1(n695), .A2(p10_mult_21_n974), .B1(p10_mult_21_n974), 
        .B2(p10_mult_21_n976), .C1(n696), .C2(p10_mult_21_n976), .ZN(
        p10_mult_21_n968) );
  NOR3_X1 U791 ( .A1(n724), .A2(n723), .A3(n725), .ZN(n696) );
  NAND2_X1 U792 ( .A1(p10_mult_21_n1138), .A2(p10_mult_21_n1139), .ZN(n726) );
  OAI21_X1 U793 ( .B1(p10_mult_21_n1138), .B2(p10_mult_21_n1139), .A(
        p10_mult_21_n1137), .ZN(n727) );
  AOI222_X1 U794 ( .A1(p10_mult_21_n926), .A2(p10_mult_21_n927), .B1(
        p10_mult_21_n926), .B2(p10_mult_21_n928), .C1(p10_mult_21_n927), .C2(
        p10_mult_21_n928), .ZN(p10_mult_21_n908) );
  OAI21_X1 U795 ( .B1(p10_mult_21_n1027), .B2(p10_mult_21_n1028), .A(
        p10_mult_21_n1026), .ZN(n729) );
  OAI21_X1 U796 ( .B1(p10_mult_21_n1143), .B2(p10_mult_21_n1142), .A(
        p10_mult_21_n1141), .ZN(n731) );
  OAI21_X1 U797 ( .B1(p10_mult_21_n1180), .B2(p10_mult_21_n1179), .A(
        p10_mult_21_n1178), .ZN(n733) );
  OAI221_X1 U798 ( .B1(n912), .B2(n902), .C1(reg4[10]), .C2(reg4[11]), .A(
        p10_mult_21_n911), .ZN(p10_mult_21_n903) );
  OAI221_X1 U799 ( .B1(n903), .B2(p10_mult_21_n1287), .C1(reg4[13]), .C2(A2[0]), .A(p10_mult_21_n863), .ZN(p10_mult_21_n1378) );
  AOI221_X1 U800 ( .B1(reg4[11]), .B2(A2[0]), .C1(n902), .C2(p10_mult_21_n1287), .A(p10_mult_21_n903), .ZN(p10_mult_21_n1391) );
  AOI221_X1 U801 ( .B1(reg4[5]), .B2(A2[0]), .C1(p10_mult_21_n1046), .C2(
        p10_mult_21_n1287), .A(p10_mult_21_n1044), .ZN(p10_mult_21_n1301) );
  XOR2_X1 U802 ( .A(p10_mult_21_n1258), .B(p10_mult_21_n1259), .Z(
        p10_mult_21_n1257) );
  XOR2_X1 U803 ( .A(p10_mult_21_n1228), .B(p10_mult_21_n1229), .Z(
        p10_mult_21_n1216) );
  NAND2_X1 U804 ( .A1(p10_mult_21_n1180), .A2(p10_mult_21_n1179), .ZN(n732) );
  NAND2_X1 U805 ( .A1(p10_mult_21_n1143), .A2(p10_mult_21_n1142), .ZN(n730) );
  AOI222_X1 U806 ( .A1(p10_mult_21_n1033), .A2(p10_mult_21_n1034), .B1(
        p10_mult_21_n1033), .B2(p10_mult_21_n1035), .C1(p10_mult_21_n1034), 
        .C2(p10_mult_21_n1035), .ZN(n698) );
  NAND2_X1 U807 ( .A1(n698), .A2(p10_mult_21_n1028), .ZN(n728) );
  AOI222_X1 U808 ( .A1(p10_mult_21_n977), .A2(p10_mult_21_n978), .B1(
        p10_mult_21_n977), .B2(p10_mult_21_n979), .C1(p10_mult_21_n978), .C2(
        p10_mult_21_n979), .ZN(p10_mult_21_n967) );
  AOI222_X1 U809 ( .A1(p10_mult_21_n922), .A2(p10_mult_21_n923), .B1(
        p10_mult_21_n922), .B2(p10_mult_21_n924), .C1(p10_mult_21_n923), .C2(
        p10_mult_21_n924), .ZN(p10_mult_21_n889) );
  AOI21_X1 U810 ( .B1(p10_mult_21_n907), .B2(p10_mult_21_n909), .A(n716), .ZN(
        n717) );
  NAND2_X1 U811 ( .A1(p10_mult_21_n885), .A2(p10_mult_21_n883), .ZN(n706) );
  NAND2_X1 U812 ( .A1(p10_mult_21_n869), .A2(p10_mult_21_n871), .ZN(n709) );
  OAI21_X1 U813 ( .B1(p10_mult_21_n863), .B2(p10_mult_21_n862), .A(
        p10_mult_21_n864), .ZN(n702) );
  AND2_X1 U814 ( .A1(n683), .A2(p10_mult_21_n907), .ZN(n714) );
  OAI221_X1 U815 ( .B1(n910), .B2(p10_mult_21_n1046), .C1(reg4[4]), .C2(
        reg4[5]), .A(p10_mult_21_n1082), .ZN(p10_mult_21_n1044) );
  XOR2_X1 U816 ( .A(p10_mult_21_n1030), .B(p10_mult_21_n1039), .Z(
        p10_mult_21_n1028) );
  AND2_X1 U817 ( .A1(n698), .A2(p10_mult_21_n1026), .ZN(n724) );
  AND2_X1 U818 ( .A1(n698), .A2(p10_mult_21_n1028), .ZN(n723) );
  OAI22_X1 U819 ( .A1(n910), .A2(n889), .B1(reg4[3]), .B2(reg4[4]), .ZN(
        p10_mult_21_n1082) );
  INV_X1 U820 ( .A(p10_mult_21_n1082), .ZN(p10_mult_21_n1021) );
  INV_X1 U821 ( .A(A2[3]), .ZN(p10_mult_21_n1121) );
  INV_X1 U822 ( .A(p10_mult_21_n1165), .ZN(p10_mult_21_n1089) );
  INV_X1 U823 ( .A(p10_mult_21_n1296), .ZN(p10_mult_21_n843) );
  OR2_X1 U824 ( .A1(p10_mult_21_n1279), .A2(p10_mult_21_n1280), .ZN(n690) );
  INV_X1 U825 ( .A(p10_mult_21_n1282), .ZN(p10_mult_21_n1281) );
  AND2_X1 U826 ( .A1(p10_mult_21_n1266), .A2(p10_mult_21_n1267), .ZN(n680) );
  AND2_X1 U827 ( .A1(p10_mult_21_n1300), .A2(p10_mult_21_n1021), .ZN(n693) );
  AND2_X1 U828 ( .A1(p10_mult_21_n1266), .A2(p10_mult_21_n1268), .ZN(n679) );
  AND2_X1 U829 ( .A1(p10_mult_21_n1268), .A2(p10_mult_21_n1267), .ZN(n678) );
  AND2_X1 U830 ( .A1(p10_mult_21_n1255), .A2(p10_mult_21_n1256), .ZN(n677) );
  AND2_X1 U831 ( .A1(p10_mult_21_n1255), .A2(p10_mult_21_n1257), .ZN(n676) );
  AND2_X1 U832 ( .A1(p10_mult_21_n1256), .A2(p10_mult_21_n1257), .ZN(n675) );
  AND2_X1 U833 ( .A1(n733), .A2(n732), .ZN(p10_mult_21_n1141) );
  AND2_X1 U834 ( .A1(n731), .A2(n730), .ZN(p10_mult_21_n1138) );
  AND2_X1 U835 ( .A1(p10_mult_21_n1028), .A2(p10_mult_21_n1026), .ZN(n725) );
  AND2_X1 U836 ( .A1(n683), .A2(p10_mult_21_n909), .ZN(n715) );
  INV_X1 U837 ( .A(p10_mult_21_n889), .ZN(n716) );
  INV_X1 U838 ( .A(n717), .ZN(n713) );
  OR3_X1 U839 ( .A1(n714), .A2(n715), .A3(n713), .ZN(n685) );
  AND3_X1 U840 ( .A1(n684), .A2(n686), .A3(n685), .ZN(n688) );
  AND3_X1 U841 ( .A1(n685), .A2(n686), .A3(n684), .ZN(n687) );
  AND2_X1 U842 ( .A1(n706), .A2(p10_mult_21_n869), .ZN(n734) );
  AND3_X1 U843 ( .A1(n711), .A2(n710), .A3(n709), .ZN(p10_mult_21_n861) );
  AND2_X1 U844 ( .A1(p10_mult_21_n861), .A2(p10_mult_21_n860), .ZN(n701) );
  INV_X1 U845 ( .A(p10_mult_21_n857), .ZN(n700) );
  INV_X1 U846 ( .A(n702), .ZN(n703) );
  CLKBUF_X1 U847 ( .A(p10_mult_21_n908), .Z(n697) );
  AOI222_X4 U848 ( .A1(p10_mult_21_n1098), .A2(p10_mult_21_n1099), .B1(
        p10_mult_21_n1098), .B2(p10_mult_21_n1100), .C1(p10_mult_21_n1099), 
        .C2(p10_mult_21_n1100), .ZN(p10_mult_21_n1034) );
  AND3_X2 U849 ( .A1(n722), .A2(n720), .A3(n721), .ZN(p10_mult_21_n927) );
  OAI221_X4 U850 ( .B1(n911), .B2(n889), .C1(reg4[2]), .C2(reg4[3]), .A(
        p10_mult_21_n1165), .ZN(p10_mult_21_n1113) );
  INV_X1 U851 ( .A(p10_mult_21_n1022), .ZN(n735) );
  INV_X2 U852 ( .A(A2[0]), .ZN(p10_mult_21_n1287) );
  AOI222_X1 U853 ( .A1(p10_mult_21_n1033), .A2(p10_mult_21_n1034), .B1(
        p10_mult_21_n1033), .B2(p10_mult_21_n1035), .C1(p10_mult_21_n1034), 
        .C2(p10_mult_21_n1035), .ZN(p10_mult_21_n1027) );
  NAND2_X1 U854 ( .A1(reg2[1]), .A2(p11_mult_21_n693), .ZN(p11_mult_21_n691)
         );
  XNOR2_X1 U855 ( .A(A1[2]), .B(reg2[1]), .ZN(p11_mult_21_n690) );
  XNOR2_X1 U856 ( .A(A1[4]), .B(reg2[1]), .ZN(p11_mult_21_n694) );
  XNOR2_X1 U857 ( .A(A1[3]), .B(reg2[1]), .ZN(p11_mult_21_n692) );
  OAI22_X1 U858 ( .A1(p11_mult_21_n709), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n710), .ZN(p11_mult_21_n405) );
  XNOR2_X1 U859 ( .A(A1[6]), .B(reg2[1]), .ZN(p11_mult_21_n696) );
  XNOR2_X1 U860 ( .A(A1[5]), .B(reg2[1]), .ZN(p11_mult_21_n695) );
  XNOR2_X1 U861 ( .A(A1[7]), .B(reg2[1]), .ZN(p11_mult_21_n697) );
  OAI22_X1 U862 ( .A1(p11_mult_21_n711), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n712), .ZN(p11_mult_21_n403) );
  OAI22_X1 U863 ( .A1(p11_mult_21_n710), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n711), .ZN(p11_mult_21_n404) );
  XNOR2_X1 U864 ( .A(A1[8]), .B(reg2[1]), .ZN(p11_mult_21_n698) );
  OAI22_X1 U865 ( .A1(p11_mult_21_n712), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n713), .ZN(p11_mult_21_n402) );
  XNOR2_X1 U866 ( .A(A1[10]), .B(reg2[1]), .ZN(p11_mult_21_n700) );
  XNOR2_X1 U867 ( .A(A1[9]), .B(reg2[1]), .ZN(p11_mult_21_n699) );
  OAI22_X1 U868 ( .A1(p11_mult_21_n713), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n714), .ZN(p11_mult_21_n401) );
  XNOR2_X1 U869 ( .A(A1[11]), .B(reg2[1]), .ZN(p11_mult_21_n701) );
  OAI22_X1 U870 ( .A1(p11_mult_21_n714), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n715), .ZN(p11_mult_21_n400) );
  XNOR2_X1 U871 ( .A(A1[12]), .B(reg2[1]), .ZN(p11_mult_21_n702) );
  OAI22_X1 U872 ( .A1(p11_mult_21_n715), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n716), .ZN(p11_mult_21_n399) );
  OAI22_X1 U873 ( .A1(p11_mult_21_n717), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n718), .ZN(p11_mult_21_n397) );
  OAI22_X1 U874 ( .A1(p11_mult_21_n716), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n717), .ZN(p11_mult_21_n398) );
  OAI22_X1 U875 ( .A1(p11_mult_21_n718), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n719), .ZN(p11_mult_21_n396) );
  NAND2_X1 U876 ( .A1(p11_mult_21_n636), .A2(p11_mult_21_n299), .ZN(
        p11_mult_21_n641) );
  NAND2_X1 U877 ( .A1(p11_mult_21_n636), .A2(p11_mult_21_n294), .ZN(
        p11_mult_21_n640) );
  OAI22_X1 U878 ( .A1(p11_mult_21_n719), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n720), .ZN(p11_mult_21_n395) );
  OAI22_X1 U879 ( .A1(p11_mult_21_n720), .A2(p11_mult_21_n707), .B1(
        p11_mult_21_n708), .B2(p11_mult_21_n722), .ZN(p11_mult_21_n231) );
  AOI21_X1 U880 ( .B1(p11_mult_21_n707), .B2(p11_mult_21_n708), .A(
        p11_mult_21_n722), .ZN(p11_mult_21_n721) );
  NAND2_X1 U881 ( .A1(p11_mult_21_n829), .A2(p11_mult_21_n277), .ZN(
        p11_mult_21_n680) );
  NAND2_X1 U882 ( .A1(p11_mult_21_n829), .A2(p11_mult_21_n268), .ZN(
        p11_mult_21_n679) );
  NAND2_X1 U883 ( .A1(p11_mult_21_n148), .A2(p11_mult_21_n245), .ZN(
        p11_mult_21_n670) );
  NAND2_X1 U884 ( .A1(p11_mult_21_n148), .A2(p11_mult_21_n234), .ZN(
        p11_mult_21_n669) );
  OAI222_X1 U885 ( .A1(p11_mult_21_n826), .A2(p11_mult_21_n827), .B1(
        p11_mult_21_n826), .B2(p11_mult_21_n828), .C1(p11_mult_21_n828), .C2(
        p11_mult_21_n827), .ZN(p11_mult_21_n659) );
  NAND2_X1 U886 ( .A1(n737), .A2(n736), .ZN(p11_mult_21_n142) );
  OAI21_X1 U887 ( .B1(p11_mult_21_n186), .B2(p11_mult_21_n193), .A(
        p11_mult_21_n143), .ZN(n737) );
  NAND2_X1 U888 ( .A1(n740), .A2(n739), .ZN(p11_mult_21_n146) );
  OAI21_X1 U889 ( .B1(p11_mult_21_n233), .B2(p11_mult_21_n222), .A(n738), .ZN(
        n740) );
  NAND3_X1 U890 ( .A1(p11_mult_21_n669), .A2(p11_mult_21_n670), .A3(
        p11_mult_21_n671), .ZN(n738) );
  NAND2_X1 U891 ( .A1(p11_mult_21_n222), .A2(p11_mult_21_n233), .ZN(n739) );
  NAND2_X1 U892 ( .A1(p11_mult_21_n186), .A2(p11_mult_21_n193), .ZN(n736) );
  XNOR2_X1 U893 ( .A(p9_mult_21_n1283), .B(p9_mult_21_n1284), .ZN(
        p9_mult_21_n1289) );
  AOI22_X1 U894 ( .A1(reg4_reg[1]), .A2(p9_mult_21_n1121), .B1(B3[3]), .B2(
        p9_mult_21_n1245), .ZN(p9_mult_21_n1296) );
  NAND2_X1 U895 ( .A1(p9_mult_21_n1244), .A2(reg4_reg[1]), .ZN(
        p9_mult_21_n1294) );
  AOI22_X1 U896 ( .A1(reg4_reg[1]), .A2(p9_mult_21_n1175), .B1(B3[2]), .B2(
        p9_mult_21_n1245), .ZN(p9_mult_21_n1295) );
  AOI22_X1 U897 ( .A1(reg4_reg[1]), .A2(p9_mult_21_n1094), .B1(B3[4]), .B2(
        p9_mult_21_n1245), .ZN(p9_mult_21_n1286) );
  OAI22_X1 U898 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1273), .B1(n772), 
        .B2(p9_mult_21_n1113), .ZN(p9_mult_21_n1277) );
  AOI22_X1 U899 ( .A1(B3[6]), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(
        p9_mult_21_n1025), .ZN(p9_mult_21_n1303) );
  AOI22_X1 U900 ( .A1(B3[5]), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(
        p9_mult_21_n1062), .ZN(p9_mult_21_n1271) );
  OAI22_X1 U901 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1272), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1273), .ZN(p9_mult_21_n1265) );
  OAI22_X1 U902 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1249), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1272), .ZN(p9_mult_21_n1253) );
  OAI22_X1 U903 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1248), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1249), .ZN(p9_mult_21_n1232) );
  OAI22_X1 U904 ( .A1(p9_mult_21_n921), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(B3[10]), .ZN(p9_mult_21_n1345) );
  OAI22_X1 U905 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1316), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1248), .ZN(p9_mult_21_n1228) );
  OAI22_X1 U906 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1331), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1316), .ZN(p9_mult_21_n1313) );
  OAI22_X1 U907 ( .A1(p9_mult_21_n897), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(B3[11]), .ZN(p9_mult_21_n1363) );
  OAI22_X1 U908 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1348), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1331), .ZN(p9_mult_21_n1206) );
  OAI22_X1 U909 ( .A1(p9_mult_21_n879), .A2(p9_mult_21_n1245), .B1(reg4_reg[1]), .B2(B3[12]), .ZN(p9_mult_21_n1374) );
  OAI22_X1 U910 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1376), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1389), .ZN(p9_mult_21_n1384) );
  OAI22_X1 U911 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1389), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1348), .ZN(p9_mult_21_n1329) );
  AOI22_X1 U912 ( .A1(B3[13]), .A2(reg4_reg[1]), .B1(p9_mult_21_n1245), .B2(
        p9_mult_21_n868), .ZN(p9_mult_21_n1167) );
  OAI22_X1 U913 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1166), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1376), .ZN(p9_mult_21_n1154) );
  OAI22_X1 U914 ( .A1(p9_mult_21_n1165), .A2(p9_mult_21_n1112), .B1(
        p9_mult_21_n1113), .B2(p9_mult_21_n1166), .ZN(p9_mult_21_n1127) );
  OAI21_X1 U915 ( .B1(reg4_reg[1]), .B2(reg4_reg[0]), .A(p9_mult_21_n1167), 
        .ZN(p9_mult_21_n1125) );
  XNOR2_X1 U916 ( .A(p9_mult_21_n926), .B(n768), .ZN(p9_mult_21_n948) );
  XNOR2_X1 U917 ( .A(p9_mult_21_n906), .B(n766), .ZN(temp4[9]) );
  OAI221_X1 U918 ( .B1(reg4_reg[3]), .B2(B3[0]), .C1(p9_mult_21_n1115), .C2(
        n770), .A(p9_mult_21_n1090), .ZN(p9_mult_21_n1297) );
  AOI22_X1 U919 ( .A1(reg4_reg[3]), .A2(n775), .B1(B3[1]), .B2(
        p9_mult_21_n1115), .ZN(p9_mult_21_n1288) );
  OAI22_X1 U920 ( .A1(p9_mult_21_n1115), .A2(p9_mult_21_n1175), .B1(B3[2]), 
        .B2(reg4_reg[3]), .ZN(p9_mult_21_n1273) );
  NOR2_X1 U921 ( .A1(p9_mult_21_n1082), .A2(n769), .ZN(p9_mult_21_n1276) );
  OAI221_X1 U922 ( .B1(p9_mult_21_n1090), .B2(p9_mult_21_n1089), .C1(
        p9_mult_21_n1090), .C2(n770), .A(reg4_reg[3]), .ZN(p9_mult_21_n1291)
         );
  OAI22_X1 U923 ( .A1(p9_mult_21_n1115), .A2(n767), .B1(B3[3]), .B2(
        reg4_reg[3]), .ZN(p9_mult_21_n1272) );
  OAI22_X1 U924 ( .A1(p9_mult_21_n1115), .A2(p9_mult_21_n1094), .B1(B3[4]), 
        .B2(reg4_reg[3]), .ZN(p9_mult_21_n1249) );
  AOI22_X1 U925 ( .A1(reg4_reg[3]), .A2(p9_mult_21_n1062), .B1(B3[5]), .B2(
        p9_mult_21_n1115), .ZN(p9_mult_21_n1248) );
  OAI22_X1 U926 ( .A1(p9_mult_21_n1025), .A2(p9_mult_21_n1115), .B1(
        reg4_reg[3]), .B2(B3[6]), .ZN(p9_mult_21_n1316) );
  OAI22_X1 U927 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1246), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1247), .ZN(p9_mult_21_n1234) );
  OAI22_X1 U928 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1247), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1299), .ZN(p9_mult_21_n1260) );
  OAI22_X1 U929 ( .A1(p9_mult_21_n983), .A2(p9_mult_21_n1115), .B1(reg4_reg[3]), .B2(B3[7]), .ZN(p9_mult_21_n1331) );
  OAI22_X1 U930 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1311), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1246), .ZN(p9_mult_21_n1226) );
  OAI22_X1 U931 ( .A1(p9_mult_21_n955), .A2(p9_mult_21_n1115), .B1(reg4_reg[3]), .B2(B3[8]), .ZN(p9_mult_21_n1348) );
  OAI22_X1 U932 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1332), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1311), .ZN(p9_mult_21_n1315) );
  OAI22_X1 U933 ( .A1(p9_mult_21_n921), .A2(p9_mult_21_n1115), .B1(reg4_reg[3]), .B2(B3[10]), .ZN(p9_mult_21_n1376) );
  AOI22_X1 U934 ( .A1(B3[9]), .A2(p9_mult_21_n1115), .B1(reg4_reg[3]), .B2(
        p9_mult_21_n935), .ZN(p9_mult_21_n1389) );
  OAI22_X1 U935 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1361), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1347), .ZN(p9_mult_21_n1344) );
  OAI22_X1 U936 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1347), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1332), .ZN(p9_mult_21_n1204) );
  AOI22_X1 U937 ( .A1(B3[11]), .A2(p9_mult_21_n1115), .B1(reg4_reg[3]), .B2(
        p9_mult_21_n897), .ZN(p9_mult_21_n1166) );
  OAI22_X1 U938 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1360), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1361), .ZN(p9_mult_21_n1354) );
  AOI22_X1 U939 ( .A1(B3[13]), .A2(reg4_reg[3]), .B1(p9_mult_21_n1115), .B2(
        p9_mult_21_n868), .ZN(p9_mult_21_n1091) );
  AOI22_X1 U940 ( .A1(B3[12]), .A2(p9_mult_21_n1115), .B1(reg4_reg[3]), .B2(
        p9_mult_21_n879), .ZN(p9_mult_21_n1112) );
  OAI22_X1 U941 ( .A1(p9_mult_21_n1082), .A2(p9_mult_21_n1043), .B1(
        p9_mult_21_n1044), .B2(p9_mult_21_n1083), .ZN(p9_mult_21_n1049) );
  AOI22_X1 U942 ( .A1(reg4_reg[5]), .A2(B3[1]), .B1(n775), .B2(
        p9_mult_21_n1046), .ZN(p9_mult_21_n1300) );
  OAI221_X1 U943 ( .B1(p9_mult_21_n1022), .B2(p9_mult_21_n1021), .C1(
        p9_mult_21_n1022), .C2(n770), .A(reg4_reg[5]), .ZN(p9_mult_21_n1275)
         );
  AOI22_X1 U944 ( .A1(reg4_reg[5]), .A2(p9_mult_21_n1175), .B1(B3[2]), .B2(
        p9_mult_21_n1046), .ZN(p9_mult_21_n1247) );
  NOR2_X1 U945 ( .A1(p9_mult_21_n1014), .A2(n769), .ZN(p9_mult_21_n1252) );
  AOI22_X1 U946 ( .A1(reg4_reg[5]), .A2(n767), .B1(B3[3]), .B2(
        p9_mult_21_n1046), .ZN(p9_mult_21_n1246) );
  OAI22_X1 U947 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1317), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1318), .ZN(p9_mult_21_n1230) );
  OAI22_X1 U948 ( .A1(p9_mult_21_n1046), .A2(p9_mult_21_n1094), .B1(B3[4]), 
        .B2(reg4_reg[5]), .ZN(p9_mult_21_n1311) );
  OAI22_X1 U949 ( .A1(p9_mult_21_n1046), .A2(p9_mult_21_n1062), .B1(B3[5]), 
        .B2(reg4_reg[5]), .ZN(p9_mult_21_n1332) );
  OAI22_X1 U950 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1346), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1333), .ZN(p9_mult_21_n1336) );
  OAI22_X1 U951 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1333), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1317), .ZN(p9_mult_21_n1314) );
  OAI22_X1 U952 ( .A1(p9_mult_21_n1046), .A2(p9_mult_21_n1025), .B1(B3[6]), 
        .B2(reg4_reg[5]), .ZN(p9_mult_21_n1347) );
  OAI22_X1 U953 ( .A1(p9_mult_21_n1046), .A2(p9_mult_21_n983), .B1(B3[7]), 
        .B2(reg4_reg[5]), .ZN(p9_mult_21_n1361) );
  OAI22_X1 U954 ( .A1(p9_mult_21_n955), .A2(p9_mult_21_n1046), .B1(reg4_reg[5]), .B2(B3[8]), .ZN(p9_mult_21_n1360) );
  OAI22_X1 U955 ( .A1(p9_mult_21_n935), .A2(reg4_reg[5]), .B1(p9_mult_21_n1046), .B2(B3[9]), .ZN(p9_mult_21_n1150) );
  OAI22_X1 U956 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1388), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1346), .ZN(p9_mult_21_n1328) );
  OAI22_X1 U957 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1375), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1388), .ZN(p9_mult_21_n1385) );
  OAI22_X1 U958 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1176), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1375), .ZN(p9_mult_21_n1153) );
  AOI22_X1 U959 ( .A1(B3[10]), .A2(reg4_reg[5]), .B1(p9_mult_21_n1046), .B2(
        p9_mult_21_n921), .ZN(p9_mult_21_n1111) );
  AOI22_X1 U960 ( .A1(B3[11]), .A2(reg4_reg[5]), .B1(p9_mult_21_n1046), .B2(
        p9_mult_21_n897), .ZN(p9_mult_21_n1084) );
  OAI22_X1 U961 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1119), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1176), .ZN(p9_mult_21_n1130) );
  AOI22_X1 U962 ( .A1(B3[12]), .A2(p9_mult_21_n1046), .B1(reg4_reg[5]), .B2(
        p9_mult_21_n879), .ZN(p9_mult_21_n1043) );
  OAI22_X1 U963 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1076), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1119), .ZN(p9_mult_21_n1072) );
  AOI22_X1 U964 ( .A1(B3[13]), .A2(reg4_reg[5]), .B1(p9_mult_21_n1046), .B2(
        p9_mult_21_n868), .ZN(p9_mult_21_n1023) );
  OAI22_X1 U965 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1042), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1076), .ZN(p9_mult_21_n1053) );
  OAI22_X1 U966 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n1015), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1042), .ZN(p9_mult_21_n1017) );
  OAI22_X1 U967 ( .A1(p9_mult_21_n1014), .A2(p9_mult_21_n984), .B1(
        p9_mult_21_n985), .B2(p9_mult_21_n1015), .ZN(p9_mult_21_n997) );
  AOI22_X1 U968 ( .A1(p9_mult_21_n1279), .A2(p9_mult_21_n1280), .B1(
        p9_mult_21_n1283), .B2(p9_mult_21_n1284), .ZN(p9_mult_21_n1282) );
  AOI222_X1 U969 ( .A1(p9_mult_21_n1235), .A2(p9_mult_21_n1236), .B1(
        p9_mult_21_n1235), .B2(p9_mult_21_n1237), .C1(p9_mult_21_n1236), .C2(
        p9_mult_21_n1237), .ZN(p9_mult_21_n1221) );
  XNOR2_X1 U970 ( .A(p9_mult_21_n1304), .B(p9_mult_21_n1212), .ZN(
        p9_mult_21_n1213) );
  NAND2_X1 U971 ( .A1(p9_mult_21_n1221), .A2(p9_mult_21_n1222), .ZN(n741) );
  NAND2_X1 U972 ( .A1(p9_mult_21_n1220), .A2(p9_mult_21_n1222), .ZN(n742) );
  NAND2_X1 U973 ( .A1(n765), .A2(p9_mult_21_n1221), .ZN(n743) );
  NOR3_X1 U974 ( .A1(n746), .A2(n745), .A3(n744), .ZN(p9_mult_21_n1195) );
  AOI222_X1 U975 ( .A1(p9_mult_21_n1255), .A2(p9_mult_21_n1256), .B1(
        p9_mult_21_n1255), .B2(p9_mult_21_n1257), .C1(p9_mult_21_n1256), .C2(
        p9_mult_21_n1257), .ZN(p9_mult_21_n1239) );
  XNOR2_X1 U976 ( .A(n748), .B(p9_mult_21_n857), .ZN(p9_mult_21_n865) );
  XNOR2_X1 U977 ( .A(p9_mult_21_n1285), .B(p9_mult_21_n1278), .ZN(
        p9_mult_21_n1280) );
  OAI211_X1 U978 ( .C1(p9_mult_21_n1089), .C2(n769), .A(p9_mult_21_n1292), .B(
        p9_mult_21_n1293), .ZN(p9_mult_21_n1290) );
  NAND2_X1 U979 ( .A1(p9_mult_21_n1289), .A2(p9_mult_21_n1291), .ZN(n747) );
  AOI222_X1 U980 ( .A1(p9_mult_21_n1258), .A2(p9_mult_21_n1261), .B1(
        p9_mult_21_n1258), .B2(p9_mult_21_n1260), .C1(p9_mult_21_n1261), .C2(
        p9_mult_21_n1260), .ZN(p9_mult_21_n1238) );
  NOR3_X1 U981 ( .A1(n751), .A2(n750), .A3(n749), .ZN(p9_mult_21_n1255) );
  XNOR2_X1 U982 ( .A(p9_mult_21_n870), .B(p9_mult_21_n869), .ZN(
        p9_mult_21_n876) );
  NAND2_X1 U983 ( .A1(p9_mult_21_n883), .A2(p9_mult_21_n885), .ZN(n756) );
  OAI21_X1 U984 ( .B1(B3[1]), .B2(p9_mult_21_n1245), .A(n769), .ZN(
        p9_mult_21_n1292) );
  OAI221_X1 U985 ( .B1(p9_mult_21_n952), .B2(p9_mult_21_n951), .C1(
        p9_mult_21_n952), .C2(n769), .A(reg4_reg[7]), .ZN(p9_mult_21_n1251) );
  XNOR2_X1 U986 ( .A(p9_mult_21_n1264), .B(p9_mult_21_n1265), .ZN(
        p9_mult_21_n1269) );
  NOR2_X1 U987 ( .A1(p9_mult_21_n911), .A2(n770), .ZN(p9_mult_21_n1337) );
  NOR2_X1 U988 ( .A1(p9_mult_21_n964), .A2(n769), .ZN(p9_mult_21_n1227) );
  OAI221_X1 U989 ( .B1(p9_mult_21_n918), .B2(p9_mult_21_n917), .C1(
        p9_mult_21_n918), .C2(n770), .A(reg4_reg[9]), .ZN(p9_mult_21_n1308) );
  OAI221_X1 U990 ( .B1(p9_mult_21_n881), .B2(p9_mult_21_n880), .C1(
        p9_mult_21_n881), .C2(n769), .A(reg4_reg[11]), .ZN(p9_mult_21_n1365)
         );
  AOI222_X1 U991 ( .A1(p9_mult_21_n1262), .A2(p9_mult_21_n1263), .B1(
        p9_mult_21_n1262), .B2(p9_mult_21_n1264), .C1(p9_mult_21_n1263), .C2(
        p9_mult_21_n1264), .ZN(p9_mult_21_n1256) );
  NOR2_X1 U992 ( .A1(p9_mult_21_n1063), .A2(n770), .ZN(p9_mult_21_n1380) );
  OAI221_X1 U993 ( .B1(p9_mult_21_n867), .B2(n769), .C1(reg4_reg[13]), .C2(
        B3[0]), .A(p9_mult_21_n863), .ZN(p9_mult_21_n1378) );
  AOI222_X1 U994 ( .A1(p9_mult_21_n886), .A2(p9_mult_21_n887), .B1(
        p9_mult_21_n886), .B2(p9_mult_21_n874), .C1(p9_mult_21_n887), .C2(
        p9_mult_21_n874), .ZN(p9_mult_21_n869) );
  NAND2_X1 U995 ( .A1(n758), .A2(p9_mult_21_n1281), .ZN(p9_mult_21_n1266) );
  NOR2_X1 U996 ( .A1(p9_mult_21_n1275), .A2(p9_mult_21_n1274), .ZN(
        p9_mult_21_n1261) );
  XNOR2_X1 U997 ( .A(p9_mult_21_n1274), .B(p9_mult_21_n1275), .ZN(
        p9_mult_21_n1264) );
  AOI21_X1 U998 ( .B1(p9_mult_21_n1300), .B2(p9_mult_21_n1021), .A(
        p9_mult_21_n1301), .ZN(p9_mult_21_n1274) );
  XNOR2_X1 U999 ( .A(p9_mult_21_n1269), .B(p9_mult_21_n1270), .ZN(
        p9_mult_21_n1268) );
  OAI22_X1 U1000 ( .A1(p9_mult_21_n987), .A2(p9_mult_21_n1121), .B1(B3[3]), 
        .B2(reg4_reg[7]), .ZN(p9_mult_21_n1333) );
  AOI22_X1 U1001 ( .A1(reg4_reg[9]), .A2(n767), .B1(B3[3]), .B2(
        p9_mult_21_n939), .ZN(p9_mult_21_n1364) );
  OAI22_X1 U1002 ( .A1(p9_mult_21_n905), .A2(B3[3]), .B1(n767), .B2(
        reg4_reg[11]), .ZN(p9_mult_21_n1149) );
  AOI22_X1 U1003 ( .A1(reg4_reg[13]), .A2(p9_mult_21_n1121), .B1(B3[3]), .B2(
        p9_mult_21_n867), .ZN(p9_mult_21_n1093) );
  AOI222_X1 U1004 ( .A1(p9_mult_21_n1276), .A2(p9_mult_21_n1277), .B1(
        p9_mult_21_n1276), .B2(p9_mult_21_n1278), .C1(p9_mult_21_n1277), .C2(
        p9_mult_21_n1278), .ZN(p9_mult_21_n1267) );
  XNOR2_X1 U1005 ( .A(p9_mult_21_n1277), .B(p9_mult_21_n1276), .ZN(
        p9_mult_21_n1285) );
  XNOR2_X1 U1006 ( .A(p9_mult_21_n1181), .B(p9_mult_21_n1182), .ZN(
        p9_mult_21_n1180) );
  NAND2_X1 U1007 ( .A1(p9_mult_21_n1179), .A2(p9_mult_21_n1180), .ZN(n761) );
  NAND2_X1 U1008 ( .A1(p9_mult_21_n1178), .A2(p9_mult_21_n1179), .ZN(n763) );
  NOR3_X1 U1009 ( .A1(n754), .A2(n753), .A3(n752), .ZN(p9_mult_21_n1220) );
  NOR3_X1 U1010 ( .A1(n754), .A2(n753), .A3(n752), .ZN(n765) );
  AOI222_X1 U1011 ( .A1(p9_mult_21_n907), .A2(p9_mult_21_n908), .B1(
        p9_mult_21_n907), .B2(p9_mult_21_n909), .C1(p9_mult_21_n908), .C2(
        p9_mult_21_n909), .ZN(n766) );
  AOI221_X1 U1012 ( .B1(reg4_reg[5]), .B2(B3[0]), .C1(p9_mult_21_n1046), .C2(
        n770), .A(p9_mult_21_n1044), .ZN(p9_mult_21_n1301) );
  NAND2_X1 U1013 ( .A1(n771), .A2(p9_mult_21_n1297), .ZN(p9_mult_21_n1283) );
  AOI22_X1 U1014 ( .A1(reg4_reg[3]), .A2(n775), .B1(B3[1]), .B2(
        p9_mult_21_n1115), .ZN(n772) );
  OAI22_X1 U1015 ( .A1(p9_mult_21_n987), .A2(n775), .B1(B3[1]), .B2(
        reg4_reg[7]), .ZN(p9_mult_21_n1318) );
  OAI22_X1 U1016 ( .A1(p9_mult_21_n939), .A2(n775), .B1(B3[1]), .B2(
        reg4_reg[9]), .ZN(p9_mult_21_n1340) );
  OAI22_X1 U1017 ( .A1(p9_mult_21_n905), .A2(B3[1]), .B1(n775), .B2(
        reg4_reg[11]), .ZN(p9_mult_21_n1390) );
  OAI22_X1 U1018 ( .A1(p9_mult_21_n867), .A2(n775), .B1(B3[1]), .B2(
        reg4_reg[13]), .ZN(p9_mult_21_n1174) );
  OAI21_X1 U1019 ( .B1(p9_mult_21_n1089), .B2(p9_mult_21_n1090), .A(
        p9_mult_21_n1091), .ZN(p9_mult_21_n1064) );
  XNOR2_X1 U1020 ( .A(p9_mult_21_n974), .B(n776), .ZN(p9_mult_21_n1002) );
  AOI222_X1 U1021 ( .A1(p9_mult_21_n974), .A2(n776), .B1(p9_mult_21_n974), 
        .B2(p9_mult_21_n976), .C1(p9_mult_21_n975), .C2(p9_mult_21_n976), .ZN(
        n774) );
  NAND2_X1 U1022 ( .A1(n780), .A2(p9_mult_21_n857), .ZN(n781) );
  XNOR2_X1 U1023 ( .A(n785), .B(n784), .ZN(temp4[13]) );
  OAI21_X1 U1024 ( .B1(p9_mult_21_n870), .B2(p9_mult_21_n871), .A(
        p9_mult_21_n869), .ZN(n778) );
  NAND2_X1 U1025 ( .A1(n782), .A2(n781), .ZN(n785) );
  OAI21_X1 U1026 ( .B1(n748), .B2(p9_mult_21_n860), .A(n777), .ZN(n782) );
  NAND3_X1 U1027 ( .A1(n779), .A2(n778), .A3(p9_mult_21_n860), .ZN(n780) );
  NAND2_X1 U1028 ( .A1(n760), .A2(p9_mult_21_n883), .ZN(n757) );
  NAND2_X1 U1029 ( .A1(p9_mult_21_n908), .A2(p9_mult_21_n907), .ZN(n786) );
  NAND2_X1 U1030 ( .A1(p9_mult_21_n908), .A2(p9_mult_21_n909), .ZN(n787) );
  NAND2_X1 U1031 ( .A1(p9_mult_21_n908), .A2(p9_mult_21_n909), .ZN(n789) );
  NAND4_X1 U1032 ( .A1(n786), .A2(n787), .A3(p9_mult_21_n890), .A4(n788), .ZN(
        n793) );
  NAND2_X1 U1033 ( .A1(p9_mult_21_n908), .A2(p9_mult_21_n907), .ZN(n790) );
  NAND3_X1 U1034 ( .A1(n814), .A2(n790), .A3(n789), .ZN(n792) );
  NOR2_X1 U1035 ( .A1(n796), .A2(n795), .ZN(n794) );
  NAND2_X1 U1036 ( .A1(n797), .A2(p9_mult_21_n890), .ZN(n800) );
  NAND2_X1 U1037 ( .A1(n794), .A2(p9_mult_21_n889), .ZN(n801) );
  NOR2_X1 U1038 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND3_X1 U1039 ( .A1(n801), .A2(n800), .A3(n799), .ZN(n755) );
  AOI222_X1 U1040 ( .A1(p9_mult_21_n967), .A2(n773), .B1(p9_mult_21_n967), 
        .B2(p9_mult_21_n969), .C1(p9_mult_21_n968), .C2(p9_mult_21_n969), .ZN(
        p9_mult_21_n927) );
  AOI222_X1 U1041 ( .A1(p9_mult_21_n974), .A2(n776), .B1(p9_mult_21_n974), 
        .B2(p9_mult_21_n976), .C1(p9_mult_21_n975), .C2(p9_mult_21_n976), .ZN(
        p9_mult_21_n968) );
  NAND2_X1 U1042 ( .A1(n774), .A2(p9_mult_21_n969), .ZN(n802) );
  NAND2_X1 U1043 ( .A1(p9_mult_21_n1138), .A2(p9_mult_21_n1139), .ZN(n803) );
  OAI21_X1 U1044 ( .B1(p9_mult_21_n1138), .B2(p9_mult_21_n1139), .A(
        p9_mult_21_n1137), .ZN(n804) );
  AOI21_X1 U1045 ( .B1(n807), .B2(n806), .A(n805), .ZN(n808) );
  NAND3_X1 U1046 ( .A1(n763), .A2(n762), .A3(n761), .ZN(n807) );
  NAND2_X1 U1047 ( .A1(p9_mult_21_n1178), .A2(p9_mult_21_n1180), .ZN(n762) );
  AOI21_X1 U1048 ( .B1(p9_mult_21_n1195), .B2(n813), .A(n812), .ZN(
        p9_mult_21_n1189) );
  OAI221_X1 U1049 ( .B1(p9_mult_21_n1395), .B2(p9_mult_21_n905), .C1(
        reg4_reg[10]), .C2(reg4_reg[11]), .A(p9_mult_21_n911), .ZN(
        p9_mult_21_n903) );
  AOI221_X1 U1050 ( .B1(reg4_reg[11]), .B2(B3[0]), .C1(p9_mult_21_n905), .C2(
        n769), .A(p9_mult_21_n903), .ZN(p9_mult_21_n1391) );
  AOI221_X1 U1051 ( .B1(reg4_reg[9]), .B2(B3[0]), .C1(p9_mult_21_n939), .C2(
        n769), .A(p9_mult_21_n937), .ZN(p9_mult_21_n1339) );
  MUX2_X1 U1052 ( .A(p9_mult_21_n842), .B(p9_mult_21_n843), .S(reg4_reg[0]), 
        .Z(p9_mult_21_n1284) );
  AOI222_X1 U1053 ( .A1(p9_mult_21_n1216), .A2(p9_mult_21_n1217), .B1(
        p9_mult_21_n1216), .B2(p9_mult_21_n1218), .C1(p9_mult_21_n1217), .C2(
        p9_mult_21_n1218), .ZN(p9_mult_21_n1215) );
  AOI222_X1 U1054 ( .A1(p9_mult_21_n1185), .A2(p9_mult_21_n1186), .B1(
        p9_mult_21_n1185), .B2(p9_mult_21_n1187), .C1(p9_mult_21_n1186), .C2(
        p9_mult_21_n1187), .ZN(p9_mult_21_n1179) );
  AOI222_X1 U1055 ( .A1(p9_mult_21_n1026), .A2(p9_mult_21_n1027), .B1(
        p9_mult_21_n1026), .B2(p9_mult_21_n1028), .C1(p9_mult_21_n1027), .C2(
        p9_mult_21_n1028), .ZN(p9_mult_21_n975) );
  AOI222_X1 U1056 ( .A1(p9_mult_21_n974), .A2(n776), .B1(p9_mult_21_n974), 
        .B2(p9_mult_21_n976), .C1(p9_mult_21_n975), .C2(p9_mult_21_n976), .ZN(
        n773) );
  NAND2_X1 U1057 ( .A1(p9_mult_21_n907), .A2(p9_mult_21_n909), .ZN(n788) );
  NAND2_X1 U1058 ( .A1(p9_mult_21_n889), .A2(p9_mult_21_n890), .ZN(n791) );
  XOR2_X1 U1059 ( .A(p9_mult_21_n895), .B(p9_mult_21_n887), .Z(p9_mult_21_n885) );
  AOI21_X1 U1060 ( .B1(p9_mult_21_n889), .B2(p9_mult_21_n890), .A(n798), .ZN(
        n799) );
  XOR2_X1 U1061 ( .A(p9_mult_21_n872), .B(p9_mult_21_n877), .Z(p9_mult_21_n871) );
  NAND2_X1 U1062 ( .A1(n759), .A2(p9_mult_21_n871), .ZN(n779) );
  OAI21_X1 U1063 ( .B1(p9_mult_21_n863), .B2(p9_mult_21_n862), .A(
        p9_mult_21_n864), .ZN(n783) );
  INV_X1 U1064 ( .A(p9_mult_21_n1082), .ZN(p9_mult_21_n1021) );
  INV_X1 U1065 ( .A(p9_mult_21_n1014), .ZN(p9_mult_21_n951) );
  INV_X1 U1066 ( .A(B3[0]), .ZN(n769) );
  INV_X1 U1067 ( .A(B3[3]), .ZN(n767) );
  INV_X1 U1068 ( .A(p9_mult_21_n1165), .ZN(p9_mult_21_n1089) );
  INV_X1 U1069 ( .A(B3[3]), .ZN(p9_mult_21_n1121) );
  INV_X1 U1070 ( .A(p9_mult_21_n1113), .ZN(p9_mult_21_n1090) );
  OR2_X1 U1071 ( .A1(p9_mult_21_n1288), .A2(p9_mult_21_n1165), .ZN(n771) );
  INV_X1 U1072 ( .A(p9_mult_21_n1296), .ZN(p9_mult_21_n843) );
  OR2_X1 U1073 ( .A1(p9_mult_21_n1280), .A2(p9_mult_21_n1279), .ZN(n758) );
  INV_X1 U1074 ( .A(p9_mult_21_n1282), .ZN(p9_mult_21_n1281) );
  AND2_X1 U1075 ( .A1(p9_mult_21_n1266), .A2(p9_mult_21_n1267), .ZN(n751) );
  AND2_X1 U1076 ( .A1(p9_mult_21_n1266), .A2(p9_mult_21_n1268), .ZN(n750) );
  AND2_X1 U1077 ( .A1(p9_mult_21_n1267), .A2(p9_mult_21_n1268), .ZN(n749) );
  INV_X1 U1078 ( .A(p9_mult_21_n1270), .ZN(p9_mult_21_n1263) );
  AND2_X1 U1079 ( .A1(p9_mult_21_n1239), .A2(p9_mult_21_n1238), .ZN(n754) );
  AND2_X1 U1080 ( .A1(p9_mult_21_n1238), .A2(p9_mult_21_n1240), .ZN(n753) );
  AND2_X1 U1081 ( .A1(p9_mult_21_n1239), .A2(p9_mult_21_n1240), .ZN(n752) );
  AND3_X1 U1082 ( .A1(n743), .A2(n742), .A3(n741), .ZN(p9_mult_21_n1214) );
  AND2_X1 U1083 ( .A1(p9_mult_21_n1213), .A2(p9_mult_21_n1214), .ZN(n746) );
  AND2_X1 U1084 ( .A1(p9_mult_21_n1213), .A2(p9_mult_21_n1215), .ZN(n745) );
  OR2_X1 U1085 ( .A1(p9_mult_21_n1196), .A2(p9_mult_21_n1197), .ZN(n813) );
  AND2_X1 U1086 ( .A1(p9_mult_21_n1196), .A2(p9_mult_21_n1197), .ZN(n812) );
  AND2_X1 U1087 ( .A1(p9_mult_21_n1189), .A2(p9_mult_21_n1190), .ZN(n809) );
  AND2_X1 U1088 ( .A1(p9_mult_21_n1189), .A2(p9_mult_21_n1188), .ZN(n810) );
  AND2_X1 U1089 ( .A1(p9_mult_21_n1190), .A2(p9_mult_21_n1188), .ZN(n811) );
  AND3_X1 U1090 ( .A1(n763), .A2(n762), .A3(n761), .ZN(n764) );
  INV_X1 U1091 ( .A(p9_mult_21_n1142), .ZN(n806) );
  INV_X1 U1092 ( .A(p9_mult_21_n1143), .ZN(n805) );
  AND2_X1 U1093 ( .A1(n788), .A2(p9_mult_21_n889), .ZN(n814) );
  AND3_X1 U1094 ( .A1(n793), .A2(n792), .A3(n791), .ZN(n760) );
  AND2_X1 U1095 ( .A1(p9_mult_21_n908), .A2(p9_mult_21_n909), .ZN(n795) );
  INV_X1 U1096 ( .A(p9_mult_21_n885), .ZN(n798) );
  AND3_X1 U1097 ( .A1(n757), .A2(n756), .A3(n755), .ZN(n759) );
  INV_X1 U1098 ( .A(p9_mult_21_n857), .ZN(n777) );
  INV_X1 U1099 ( .A(n783), .ZN(n784) );
  AOI222_X4 U1100 ( .A1(p9_mult_21_n926), .A2(n768), .B1(p9_mult_21_n926), 
        .B2(p9_mult_21_n928), .C1(p9_mult_21_n927), .C2(p9_mult_21_n928), .ZN(
        p9_mult_21_n908) );
  OAI22_X2 U1101 ( .A1(p9_mult_21_n1394), .A2(p9_mult_21_n1245), .B1(
        reg4_reg[1]), .B2(reg4_reg[2]), .ZN(p9_mult_21_n1165) );
  OAI221_X4 U1102 ( .B1(p9_mult_21_n1394), .B2(p9_mult_21_n1115), .C1(
        reg4_reg[2]), .C2(reg4_reg[3]), .A(p9_mult_21_n1165), .ZN(
        p9_mult_21_n1113) );
  OAI22_X2 U1103 ( .A1(p9_mult_21_n1370), .A2(p9_mult_21_n1115), .B1(
        reg4_reg[3]), .B2(reg4_reg[4]), .ZN(p9_mult_21_n1082) );
  AOI222_X1 U1104 ( .A1(p9_mult_21_n1033), .A2(p9_mult_21_n1034), .B1(
        p9_mult_21_n1033), .B2(p9_mult_21_n1035), .C1(p9_mult_21_n1034), .C2(
        p9_mult_21_n1035), .ZN(p9_mult_21_n1027) );
  AOI222_X4 U1105 ( .A1(p9_mult_21_n1026), .A2(p9_mult_21_n1027), .B1(
        p9_mult_21_n1026), .B2(p9_mult_21_n1028), .C1(p9_mult_21_n1027), .C2(
        p9_mult_21_n1028), .ZN(n776) );
  AND2_X2 U1106 ( .A1(n804), .A2(n803), .ZN(p9_mult_21_n1100) );
  AOI222_X2 U1107 ( .A1(p9_mult_21_n1098), .A2(p9_mult_21_n1099), .B1(
        p9_mult_21_n1098), .B2(p9_mult_21_n1100), .C1(p9_mult_21_n1099), .C2(
        p9_mult_21_n1100), .ZN(p9_mult_21_n1034) );
  AOI222_X1 U1108 ( .A1(p9_mult_21_n869), .A2(p9_mult_21_n870), .B1(
        p9_mult_21_n869), .B2(p9_mult_21_n871), .C1(n759), .C2(p9_mult_21_n871), .ZN(n748) );
  NOR3_X2 U1109 ( .A1(n809), .A2(n810), .A3(n811), .ZN(p9_mult_21_n1178) );
  AND3_X2 U1110 ( .A1(n757), .A2(n756), .A3(n755), .ZN(p9_mult_21_n870) );
  AOI21_X1 U1111 ( .B1(n764), .B2(p9_mult_21_n1142), .A(n808), .ZN(
        p9_mult_21_n1138) );
  OAI22_X2 U1112 ( .A1(p9_mult_21_n1393), .A2(p9_mult_21_n1046), .B1(
        reg4_reg[5]), .B2(reg4_reg[6]), .ZN(p9_mult_21_n1014) );
  XNOR2_X1 U1113 ( .A(B2[2]), .B(reg3_reg[3]), .ZN(p8_mult_21_n708) );
  XNOR2_X1 U1114 ( .A(B2[1]), .B(reg3_reg[3]), .ZN(p8_mult_21_n707) );
  XNOR2_X1 U1115 ( .A(reg3_reg[3]), .B(B2[0]), .ZN(p8_mult_21_n704) );
  NOR2_X1 U1116 ( .A1(p8_mult_21_n721), .A2(p8_mult_21_n722), .ZN(
        p8_mult_21_n393) );
  XNOR2_X1 U1117 ( .A(B2[4]), .B(reg3_reg[3]), .ZN(p8_mult_21_n710) );
  XNOR2_X1 U1118 ( .A(B2[3]), .B(reg3_reg[3]), .ZN(p8_mult_21_n709) );
  XNOR2_X1 U1119 ( .A(B2[5]), .B(reg3_reg[3]), .ZN(p8_mult_21_n711) );
  OAI22_X1 U1120 ( .A1(p8_mult_21_n726), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n727), .ZN(p8_mult_21_n390) );
  XNOR2_X1 U1121 ( .A(B2[6]), .B(reg3_reg[3]), .ZN(p8_mult_21_n712) );
  OAI22_X1 U1122 ( .A1(p8_mult_21_n727), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n728), .ZN(p8_mult_21_n389) );
  XNOR2_X1 U1123 ( .A(B2[7]), .B(reg3_reg[3]), .ZN(p8_mult_21_n713) );
  XNOR2_X1 U1124 ( .A(B2[8]), .B(reg3_reg[3]), .ZN(p8_mult_21_n714) );
  OAI22_X1 U1125 ( .A1(p8_mult_21_n728), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n729), .ZN(p8_mult_21_n388) );
  XNOR2_X1 U1126 ( .A(B2[10]), .B(reg3_reg[3]), .ZN(p8_mult_21_n716) );
  XNOR2_X1 U1127 ( .A(B2[9]), .B(reg3_reg[3]), .ZN(p8_mult_21_n715) );
  OAI22_X1 U1128 ( .A1(p8_mult_21_n730), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n731), .ZN(p8_mult_21_n386) );
  OAI22_X1 U1129 ( .A1(p8_mult_21_n729), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n730), .ZN(p8_mult_21_n387) );
  XNOR2_X1 U1130 ( .A(B2[11]), .B(reg3_reg[3]), .ZN(p8_mult_21_n717) );
  OAI22_X1 U1131 ( .A1(p8_mult_21_n732), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n733), .ZN(p8_mult_21_n384) );
  XNOR2_X1 U1132 ( .A(B2[12]), .B(reg3_reg[3]), .ZN(p8_mult_21_n718) );
  OAI22_X1 U1133 ( .A1(p8_mult_21_n731), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n732), .ZN(p8_mult_21_n385) );
  NAND2_X1 U1134 ( .A1(p8_mult_21_n636), .A2(p8_mult_21_n299), .ZN(
        p8_mult_21_n641) );
  XNOR2_X1 U1135 ( .A(B2[13]), .B(reg3_reg[3]), .ZN(p8_mult_21_n720) );
  OAI22_X1 U1136 ( .A1(p8_mult_21_n733), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n734), .ZN(p8_mult_21_n817) );
  OAI22_X1 U1137 ( .A1(p8_mult_21_n734), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n735), .ZN(p8_mult_21_n382) );
  OAI22_X1 U1138 ( .A1(p8_mult_21_n735), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n736), .ZN(p8_mult_21_n381) );
  OAI22_X1 U1139 ( .A1(p8_mult_21_n736), .A2(p8_mult_21_n724), .B1(
        p8_mult_21_n722), .B2(p8_mult_21_n738), .ZN(p8_mult_21_n209) );
  AOI21_X1 U1140 ( .B1(p8_mult_21_n724), .B2(p8_mult_21_n722), .A(
        p8_mult_21_n738), .ZN(p8_mult_21_n737) );
  OAI22_X1 U1141 ( .A1(p8_mult_21_n704), .A2(p8_mult_21_n705), .B1(
        p8_mult_21_n706), .B2(p8_mult_21_n707), .ZN(p8_mult_21_n406) );
  NOR2_X1 U1142 ( .A1(p8_mult_21_n832), .A2(p8_mult_21_n681), .ZN(
        p8_mult_21_n644) );
  OAI222_X1 U1143 ( .A1(p8_mult_21_n824), .A2(p8_mult_21_n825), .B1(
        p8_mult_21_n824), .B2(p8_mult_21_n826), .C1(p8_mult_21_n826), .C2(
        p8_mult_21_n825), .ZN(p8_mult_21_n657) );
  NAND2_X1 U1144 ( .A1(n816), .A2(n815), .ZN(p8_mult_21_n142) );
  OAI21_X1 U1145 ( .B1(p8_mult_21_n186), .B2(p8_mult_21_n193), .A(
        p8_mult_21_n143), .ZN(n816) );
  NAND2_X1 U1146 ( .A1(n818), .A2(n817), .ZN(p8_mult_21_n146) );
  OAI21_X1 U1147 ( .B1(p8_mult_21_n233), .B2(p8_mult_21_n222), .A(
        p8_mult_21_n147), .ZN(n818) );
  NAND2_X1 U1148 ( .A1(n820), .A2(n819), .ZN(p8_mult_21_n147) );
  OAI21_X1 U1149 ( .B1(p8_mult_21_n245), .B2(p8_mult_21_n234), .A(
        p8_mult_21_n148), .ZN(n820) );
  NAND2_X1 U1150 ( .A1(p8_mult_21_n234), .A2(p8_mult_21_n245), .ZN(n819) );
  NAND2_X1 U1151 ( .A1(p8_mult_21_n222), .A2(p8_mult_21_n233), .ZN(n817) );
  NAND2_X1 U1152 ( .A1(p8_mult_21_n186), .A2(p8_mult_21_n193), .ZN(n815) );
  AOI222_X1 U1153 ( .A1(p7_mult_21_n1226), .A2(p7_mult_21_n1227), .B1(
        p7_mult_21_n1226), .B2(p7_mult_21_n1228), .C1(p7_mult_21_n1227), .C2(
        p7_mult_21_n1228), .ZN(p7_mult_21_n1215) );
  AOI222_X1 U1154 ( .A1(p7_mult_21_n1215), .A2(p7_mult_21_n1216), .B1(
        p7_mult_21_n1215), .B2(p7_mult_21_n1217), .C1(p7_mult_21_n1216), .C2(
        p7_mult_21_n1217), .ZN(p7_mult_21_n1214) );
  AOI222_X1 U1155 ( .A1(p7_mult_21_n1239), .A2(p7_mult_21_n1240), .B1(
        p7_mult_21_n1239), .B2(p7_mult_21_n1241), .C1(p7_mult_21_n1240), .C2(
        p7_mult_21_n1241), .ZN(p7_mult_21_n1229) );
  AOI222_X1 U1156 ( .A1(p7_mult_21_n1229), .A2(p7_mult_21_n1230), .B1(
        p7_mult_21_n1229), .B2(p7_mult_21_n1231), .C1(p7_mult_21_n1230), .C2(
        p7_mult_21_n1231), .ZN(p7_mult_21_n1228) );
  AOI222_X1 U1157 ( .A1(p7_mult_21_n1212), .A2(p7_mult_21_n1213), .B1(
        p7_mult_21_n1212), .B2(p7_mult_21_n1214), .C1(p7_mult_21_n1213), .C2(
        p7_mult_21_n1214), .ZN(p7_mult_21_n1193) );
  XNOR2_X1 U1158 ( .A(p7_mult_21_n932), .B(p7_mult_21_n933), .ZN(
        p7_mult_21_n954) );
  XNOR2_X1 U1159 ( .A(p7_mult_21_n865), .B(p7_mult_21_n869), .ZN(temp2[12]) );
  AOI22_X1 U1160 ( .A1(p7_mult_21_n1253), .A2(p7_mult_21_n1252), .B1(
        p7_mult_21_n1256), .B2(p7_mult_21_n1257), .ZN(p7_mult_21_n1255) );
  AOI22_X1 U1161 ( .A1(p7_mult_21_n1133), .A2(reg2_reg[1]), .B1(
        p7_mult_21_n1261), .B2(B1[3]), .ZN(p7_mult_21_n1273) );
  AOI22_X1 U1162 ( .A1(reg2_reg[1]), .A2(B1[4]), .B1(n841), .B2(
        p7_mult_21_n1261), .ZN(p7_mult_21_n1262) );
  AOI22_X1 U1163 ( .A1(reg2_reg[1]), .A2(p7_mult_21_n1180), .B1(B1[2]), .B2(
        p7_mult_21_n1261), .ZN(p7_mult_21_n1272) );
  AOI22_X1 U1164 ( .A1(B1[5]), .A2(reg2_reg[1]), .B1(p7_mult_21_n1261), .B2(
        p7_mult_21_n1068), .ZN(p7_mult_21_n1288) );
  AOI22_X1 U1165 ( .A1(B1[10]), .A2(reg2_reg[1]), .B1(p7_mult_21_n1261), .B2(
        p7_mult_21_n924), .ZN(p7_mult_21_n1350) );
  OAI22_X1 U1166 ( .A1(p7_mult_21_n885), .A2(p7_mult_21_n1261), .B1(
        reg2_reg[1]), .B2(B1[12]), .ZN(p7_mult_21_n1381) );
  AOI22_X1 U1167 ( .A1(B1[11]), .A2(reg2_reg[1]), .B1(p7_mult_21_n1261), .B2(
        p7_mult_21_n904), .ZN(p7_mult_21_n1370) );
  OAI22_X1 U1168 ( .A1(p7_mult_21_n877), .A2(p7_mult_21_n1261), .B1(
        reg2_reg[1]), .B2(B1[13]), .ZN(p7_mult_21_n1172) );
  OAI21_X1 U1169 ( .B1(reg2_reg[1]), .B2(reg2_reg[0]), .A(p7_mult_21_n1171), 
        .ZN(p7_mult_21_n1137) );
  XNOR2_X1 U1170 ( .A(p7_mult_21_n1257), .B(p7_mult_21_n1256), .ZN(
        p7_mult_21_n1266) );
  AOI222_X1 U1171 ( .A1(p7_mult_21_n1266), .A2(p7_mult_21_n1267), .B1(
        p7_mult_21_n1266), .B2(p7_mult_21_n1268), .C1(p7_mult_21_n1267), .C2(
        p7_mult_21_n1268), .ZN(p7_mult_21_n1252) );
  AOI222_X1 U1172 ( .A1(p7_mult_21_n1243), .A2(p7_mult_21_n1242), .B1(
        p7_mult_21_n1242), .B2(p7_mult_21_n1244), .C1(p7_mult_21_n1244), .C2(
        p7_mult_21_n1243), .ZN(p7_mult_21_n1241) );
  AOI22_X1 U1173 ( .A1(reg2_reg[3]), .A2(n829), .B1(B1[3]), .B2(
        p7_mult_21_n1126), .ZN(p7_mult_21_n1287) );
  AOI22_X1 U1174 ( .A1(reg2_reg[5]), .A2(n829), .B1(B1[3]), .B2(
        p7_mult_21_n1053), .ZN(p7_mult_21_n1305) );
  OAI22_X1 U1175 ( .A1(p7_mult_21_n992), .A2(n829), .B1(B1[3]), .B2(
        reg2_reg[7]), .ZN(p7_mult_21_n1343) );
  AOI22_X1 U1176 ( .A1(reg2_reg[9]), .A2(n829), .B1(B1[3]), .B2(
        p7_mult_21_n945), .ZN(p7_mult_21_n1372) );
  OAI22_X1 U1177 ( .A1(p7_mult_21_n911), .A2(B1[3]), .B1(n829), .B2(
        reg2_reg[11]), .ZN(p7_mult_21_n1155) );
  AOI22_X1 U1178 ( .A1(reg2_reg[13]), .A2(n829), .B1(B1[3]), .B2(
        p7_mult_21_n876), .ZN(p7_mult_21_n1099) );
  OAI221_X1 U1179 ( .B1(reg2_reg[3]), .B2(B1[0]), .C1(p7_mult_21_n1126), .C2(
        n831), .A(p7_mult_21_n1096), .ZN(p7_mult_21_n1274) );
  OAI221_X1 U1180 ( .B1(reg2_reg[5]), .B2(B1[0]), .C1(p7_mult_21_n1053), .C2(
        n830), .A(p7_mult_21_n1029), .ZN(p7_mult_21_n1285) );
  OAI21_X1 U1181 ( .B1(B1[1]), .B2(p7_mult_21_n1261), .A(n831), .ZN(
        p7_mult_21_n1269) );
  NOR2_X1 U1182 ( .A1(p7_mult_21_n1089), .A2(n830), .ZN(p7_mult_21_n1245) );
  OAI21_X1 U1183 ( .B1(p7_mult_21_n1265), .B2(p7_mult_21_n1169), .A(
        p7_mult_21_n1274), .ZN(p7_mult_21_n1256) );
  OAI221_X1 U1184 ( .B1(p7_mult_21_n1096), .B2(p7_mult_21_n1095), .C1(
        p7_mult_21_n1096), .C2(n830), .A(reg2_reg[3]), .ZN(p7_mult_21_n1268)
         );
  OAI211_X1 U1185 ( .C1(p7_mult_21_n1095), .C2(n831), .A(p7_mult_21_n1269), 
        .B(p7_mult_21_n1270), .ZN(p7_mult_21_n1267) );
  NOR2_X1 U1186 ( .A1(p7_mult_21_n1022), .A2(n830), .ZN(p7_mult_21_n1281) );
  OAI221_X1 U1187 ( .B1(p7_mult_21_n970), .B2(n830), .C1(p7_mult_21_n919), 
        .C2(p7_mult_21_n1331), .A(reg2_reg[9]), .ZN(p7_mult_21_n1312) );
  NOR2_X1 U1188 ( .A1(p7_mult_21_n970), .A2(n831), .ZN(p7_mult_21_n1294) );
  NOR2_X1 U1189 ( .A1(p7_mult_21_n914), .A2(n831), .ZN(p7_mult_21_n1317) );
  OAI221_X1 U1190 ( .B1(p7_mult_21_n887), .B2(p7_mult_21_n886), .C1(
        p7_mult_21_n887), .C2(n830), .A(reg2_reg[11]), .ZN(p7_mult_21_n1373)
         );
  NOR2_X1 U1191 ( .A1(p7_mult_21_n883), .A2(n830), .ZN(p7_mult_21_n1387) );
  XNOR2_X1 U1192 ( .A(p7_mult_21_n1072), .B(p7_mult_21_n1042), .ZN(temp2[3])
         );
  XNOR2_X1 U1193 ( .A(p7_mult_21_n1146), .B(n843), .ZN(temp2[1]) );
  XNOR2_X1 U1194 ( .A(p7_mult_21_n895), .B(p7_mult_21_n896), .ZN(
        p7_mult_21_n912) );
  XNOR2_X1 U1195 ( .A(p7_mult_21_n1258), .B(p7_mult_21_n1247), .ZN(
        p7_mult_21_n1253) );
  XNOR2_X1 U1196 ( .A(p7_mult_21_n1114), .B(p7_mult_21_n1106), .ZN(
        p7_mult_21_n1075) );
  AOI222_X1 U1197 ( .A1(p7_mult_21_n1111), .A2(p7_mult_21_n1112), .B1(
        p7_mult_21_n1111), .B2(p7_mult_21_n1113), .C1(p7_mult_21_n1112), .C2(
        p7_mult_21_n1113), .ZN(p7_mult_21_n1073) );
  NAND2_X1 U1198 ( .A1(p7_mult_21_n1254), .A2(n822), .ZN(p7_mult_21_n1242) );
  NAND2_X1 U1199 ( .A1(p7_mult_21_n1073), .A2(p7_mult_21_n1075), .ZN(n824) );
  AOI222_X1 U1200 ( .A1(p7_mult_21_n1245), .A2(p7_mult_21_n1246), .B1(
        p7_mult_21_n1245), .B2(p7_mult_21_n1247), .C1(p7_mult_21_n1247), .C2(
        p7_mult_21_n1246), .ZN(p7_mult_21_n1244) );
  AOI22_X1 U1201 ( .A1(reg2_reg[0]), .A2(p7_mult_21_n1288), .B1(
        p7_mult_21_n1289), .B2(p7_mult_21_n1262), .ZN(p7_mult_21_n1248) );
  OAI21_X1 U1202 ( .B1(p7_mult_21_n1280), .B2(p7_mult_21_n1089), .A(
        p7_mult_21_n1285), .ZN(p7_mult_21_n1278) );
  XNOR2_X1 U1203 ( .A(p7_mult_21_n1277), .B(p7_mult_21_n1278), .ZN(
        p7_mult_21_n1251) );
  OAI22_X1 U1204 ( .A1(p7_mult_21_n1089), .A2(p7_mult_21_n1279), .B1(
        p7_mult_21_n1051), .B2(p7_mult_21_n1280), .ZN(p7_mult_21_n1234) );
  AOI22_X1 U1205 ( .A1(reg2_reg[5]), .A2(n837), .B1(B1[1]), .B2(
        p7_mult_21_n1053), .ZN(p7_mult_21_n1280) );
  XNOR2_X1 U1206 ( .A(p7_mult_21_n1250), .B(p7_mult_21_n1251), .ZN(n826) );
  XNOR2_X1 U1207 ( .A(p7_mult_21_n1248), .B(n826), .ZN(p7_mult_21_n1243) );
  AOI222_X1 U1208 ( .A1(p7_mult_21_n1232), .A2(p7_mult_21_n1233), .B1(
        p7_mult_21_n1232), .B2(p7_mult_21_n1234), .C1(p7_mult_21_n1233), .C2(
        p7_mult_21_n1234), .ZN(p7_mult_21_n1231) );
  AOI22_X1 U1209 ( .A1(reg2_reg[3]), .A2(n836), .B1(B1[1]), .B2(
        p7_mult_21_n1126), .ZN(p7_mult_21_n1265) );
  OAI22_X1 U1210 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1264), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1265), .ZN(p7_mult_21_n1246) );
  OAI22_X1 U1211 ( .A1(p7_mult_21_n1126), .A2(p7_mult_21_n1180), .B1(B1[2]), 
        .B2(reg2_reg[3]), .ZN(p7_mult_21_n1264) );
  AOI22_X1 U1212 ( .A1(reg2_reg[3]), .A2(n841), .B1(B1[4]), .B2(
        p7_mult_21_n1126), .ZN(p7_mult_21_n1308) );
  OAI22_X1 U1213 ( .A1(p7_mult_21_n1053), .A2(n841), .B1(B1[4]), .B2(
        reg2_reg[5]), .ZN(p7_mult_21_n1335) );
  OAI22_X1 U1214 ( .A1(p7_mult_21_n992), .A2(n841), .B1(B1[4]), .B2(
        reg2_reg[7]), .ZN(p7_mult_21_n1351) );
  OAI22_X1 U1215 ( .A1(p7_mult_21_n945), .A2(n841), .B1(B1[4]), .B2(
        reg2_reg[9]), .ZN(p7_mult_21_n1377) );
  AOI22_X1 U1216 ( .A1(reg2_reg[11]), .A2(B1[4]), .B1(n841), .B2(
        p7_mult_21_n911), .ZN(p7_mult_21_n1128) );
  OAI22_X1 U1217 ( .A1(p7_mult_21_n876), .A2(B1[4]), .B1(n841), .B2(
        reg2_reg[13]), .ZN(p7_mult_21_n1067) );
  XNOR2_X1 U1218 ( .A(p7_mult_21_n1246), .B(p7_mult_21_n1245), .ZN(
        p7_mult_21_n1258) );
  OAI22_X1 U1219 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1287), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1264), .ZN(p7_mult_21_n1286) );
  OAI22_X1 U1220 ( .A1(B1[1]), .A2(p7_mult_21_n1271), .B1(p7_mult_21_n1272), 
        .B2(p7_mult_21_n1260), .ZN(p7_mult_21_n1270) );
  OAI22_X1 U1221 ( .A1(p7_mult_21_n992), .A2(n835), .B1(B1[2]), .B2(
        reg2_reg[7]), .ZN(p7_mult_21_n1337) );
  AOI22_X1 U1222 ( .A1(reg2_reg[5]), .A2(n835), .B1(B1[2]), .B2(
        p7_mult_21_n1053), .ZN(p7_mult_21_n1279) );
  AOI22_X1 U1223 ( .A1(reg2_reg[9]), .A2(B1[2]), .B1(n835), .B2(
        p7_mult_21_n945), .ZN(p7_mult_21_n1356) );
  AOI22_X1 U1224 ( .A1(reg2_reg[11]), .A2(B1[2]), .B1(n835), .B2(
        p7_mult_21_n911), .ZN(p7_mult_21_n1379) );
  OAI22_X1 U1225 ( .A1(p7_mult_21_n876), .A2(n835), .B1(B1[2]), .B2(
        reg2_reg[13]), .ZN(p7_mult_21_n1132) );
  AOI222_X1 U1226 ( .A1(p7_mult_21_n1248), .A2(p7_mult_21_n1250), .B1(
        p7_mult_21_n1248), .B2(p7_mult_21_n1251), .C1(p7_mult_21_n1250), .C2(
        p7_mult_21_n1251), .ZN(p7_mult_21_n1239) );
  OAI221_X1 U1227 ( .B1(p7_mult_21_n992), .B2(n831), .C1(reg2_reg[7]), .C2(
        B1[0]), .A(p7_mult_21_n958), .ZN(p7_mult_21_n1339) );
  OAI221_X1 U1228 ( .B1(p7_mult_21_n876), .B2(n831), .C1(reg2_reg[13]), .C2(
        B1[0]), .A(p7_mult_21_n867), .ZN(p7_mult_21_n1385) );
  AOI221_X1 U1229 ( .B1(p7_mult_21_n874), .B2(p7_mult_21_n883), .C1(
        p7_mult_21_n874), .C2(B1[0]), .A(p7_mult_21_n876), .ZN(
        p7_mult_21_n1177) );
  AOI221_X1 U1230 ( .B1(p7_mult_21_n990), .B2(p7_mult_21_n1022), .C1(
        p7_mult_21_n990), .C2(B1[0]), .A(p7_mult_21_n992), .ZN(
        p7_mult_21_n1302) );
  XNOR2_X1 U1231 ( .A(p7_mult_21_n980), .B(p7_mult_21_n979), .ZN(
        p7_mult_21_n1009) );
  XNOR2_X1 U1232 ( .A(p7_mult_21_n1221), .B(p7_mult_21_n1218), .ZN(
        p7_mult_21_n1290) );
  NOR2_X1 U1233 ( .A1(B1[2]), .A2(p7_mult_21_n1261), .ZN(p7_mult_21_n846) );
  NOR2_X1 U1234 ( .A1(B1[3]), .A2(p7_mult_21_n1261), .ZN(p7_mult_21_n844) );
  NAND2_X1 U1235 ( .A1(n833), .A2(n834), .ZN(p7_mult_21_n1257) );
  NAND2_X1 U1236 ( .A1(p7_mult_21_n847), .A2(reg2_reg[0]), .ZN(n833) );
  NAND2_X1 U1237 ( .A1(p7_mult_21_n846), .A2(p7_mult_21_n1260), .ZN(n834) );
  AOI222_X1 U1238 ( .A1(p7_mult_21_n895), .A2(p7_mult_21_n896), .B1(
        p7_mult_21_n895), .B2(p7_mult_21_n897), .C1(p7_mult_21_n896), .C2(
        p7_mult_21_n897), .ZN(p7_mult_21_n890) );
  OAI22_X1 U1239 ( .A1(p7_mult_21_n992), .A2(n836), .B1(B1[1]), .B2(
        reg2_reg[7]), .ZN(p7_mult_21_n1338) );
  AOI22_X1 U1240 ( .A1(reg2_reg[9]), .A2(B1[1]), .B1(n837), .B2(
        p7_mult_21_n945), .ZN(p7_mult_21_n1332) );
  OAI22_X1 U1241 ( .A1(p7_mult_21_n911), .A2(B1[1]), .B1(n836), .B2(
        reg2_reg[11]), .ZN(p7_mult_21_n1397) );
  OAI22_X1 U1242 ( .A1(p7_mult_21_n876), .A2(n837), .B1(B1[1]), .B2(
        reg2_reg[13]), .ZN(p7_mult_21_n1179) );
  OAI22_X1 U1243 ( .A1(p7_mult_21_n1032), .A2(p7_mult_21_n1126), .B1(
        reg2_reg[3]), .B2(B1[6]), .ZN(p7_mult_21_n1336) );
  AOI22_X1 U1244 ( .A1(reg2_reg[5]), .A2(B1[6]), .B1(p7_mult_21_n1032), .B2(
        p7_mult_21_n1053), .ZN(p7_mult_21_n1353) );
  OAI22_X1 U1245 ( .A1(p7_mult_21_n992), .A2(p7_mult_21_n1032), .B1(B1[6]), 
        .B2(reg2_reg[7]), .ZN(p7_mult_21_n1382) );
  OAI22_X1 U1246 ( .A1(p7_mult_21_n945), .A2(p7_mult_21_n1032), .B1(B1[6]), 
        .B2(reg2_reg[9]), .ZN(p7_mult_21_n1130) );
  OAI22_X1 U1247 ( .A1(p7_mult_21_n911), .A2(p7_mult_21_n1032), .B1(B1[6]), 
        .B2(reg2_reg[11]), .ZN(p7_mult_21_n1054) );
  AOI22_X1 U1248 ( .A1(reg2_reg[13]), .A2(B1[6]), .B1(p7_mult_21_n1032), .B2(
        p7_mult_21_n876), .ZN(p7_mult_21_n987) );
  AOI222_X1 U1249 ( .A1(p7_mult_21_n1036), .A2(p7_mult_21_n1037), .B1(
        p7_mult_21_n1036), .B2(p7_mult_21_n1038), .C1(p7_mult_21_n1037), .C2(
        p7_mult_21_n1038), .ZN(p7_mult_21_n979) );
  OAI22_X1 U1250 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1307), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1308), .ZN(p7_mult_21_n1299) );
  OAI22_X1 U1251 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1344), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1336), .ZN(p7_mult_21_n1318) );
  OAI22_X1 U1252 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1170), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1383), .ZN(p7_mult_21_n1159) );
  OAI22_X1 U1253 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1123), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1170), .ZN(p7_mult_21_n1139) );
  OAI21_X1 U1254 ( .B1(p7_mult_21_n1123), .B2(p7_mult_21_n1124), .A(
        p7_mult_21_n1125), .ZN(p7_mult_21_n1071) );
  OAI22_X1 U1255 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1383), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1396), .ZN(p7_mult_21_n1391) );
  OAI22_X1 U1256 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1336), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1307), .ZN(p7_mult_21_n1295) );
  OAI22_X1 U1257 ( .A1(p7_mult_21_n1169), .A2(p7_mult_21_n1308), .B1(
        p7_mult_21_n1124), .B2(p7_mult_21_n1287), .ZN(p7_mult_21_n1283) );
  AOI22_X1 U1258 ( .A1(p7_mult_21_n1095), .A2(p7_mult_21_n1354), .B1(
        p7_mult_21_n1096), .B2(p7_mult_21_n1355), .ZN(p7_mult_21_n1324) );
  NAND2_X1 U1259 ( .A1(p7_mult_21_n1097), .A2(p7_mult_21_n1095), .ZN(
        p7_mult_21_n1125) );
  OAI21_X1 U1260 ( .B1(p7_mult_21_n1095), .B2(p7_mult_21_n1096), .A(
        p7_mult_21_n1097), .ZN(p7_mult_21_n1069) );
  AOI22_X1 U1261 ( .A1(p7_mult_21_n1095), .A2(p7_mult_21_n1395), .B1(
        p7_mult_21_n1096), .B2(p7_mult_21_n1354), .ZN(p7_mult_21_n1207) );
  XNOR2_X1 U1262 ( .A(p7_mult_21_n1283), .B(p7_mult_21_n1284), .ZN(n842) );
  XNOR2_X1 U1263 ( .A(p7_mult_21_n1281), .B(n842), .ZN(p7_mult_21_n1233) );
  AOI222_X1 U1264 ( .A1(p7_mult_21_n1183), .A2(p7_mult_21_n1184), .B1(
        p7_mult_21_n1183), .B2(p7_mult_21_n1185), .C1(p7_mult_21_n1184), .C2(
        p7_mult_21_n1185), .ZN(n844) );
  XNOR2_X1 U1265 ( .A(p7_mult_21_n1234), .B(p7_mult_21_n1232), .ZN(n845) );
  XNOR2_X1 U1266 ( .A(p7_mult_21_n1233), .B(n845), .ZN(p7_mult_21_n1240) );
  AOI22_X1 U1267 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1353), .B1(
        p7_mult_21_n1029), .B2(p7_mult_21_n1342), .ZN(p7_mult_21_n1322) );
  AOI22_X1 U1268 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1156), .B1(
        p7_mult_21_n1029), .B2(p7_mult_21_n1368), .ZN(p7_mult_21_n1161) );
  AOI22_X1 U1269 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1122), .B1(
        p7_mult_21_n1029), .B2(p7_mult_21_n1156), .ZN(p7_mult_21_n1135) );
  NAND2_X1 U1270 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1030), .ZN(
        p7_mult_21_n1052) );
  OAI21_X1 U1271 ( .B1(p7_mult_21_n1028), .B2(p7_mult_21_n1029), .A(
        p7_mult_21_n1030), .ZN(p7_mult_21_n998) );
  AOI22_X1 U1272 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1121), .B1(
        p7_mult_21_n1029), .B2(p7_mult_21_n1122), .ZN(p7_mult_21_n1081) );
  AOI22_X1 U1273 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1368), .B1(
        p7_mult_21_n1029), .B2(p7_mult_21_n1369), .ZN(p7_mult_21_n1361) );
  AOI22_X1 U1274 ( .A1(p7_mult_21_n1028), .A2(p7_mult_21_n1369), .B1(
        p7_mult_21_n1029), .B2(p7_mult_21_n1353), .ZN(p7_mult_21_n1348) );
  XNOR2_X1 U1275 ( .A(n846), .B(n847), .ZN(temp2[13]) );
  XOR2_X1 U1276 ( .A(n850), .B(n849), .Z(n847) );
  NAND2_X1 U1277 ( .A1(p7_mult_21_n865), .A2(p7_mult_21_n860), .ZN(n848) );
  NAND2_X1 U1278 ( .A1(n852), .A2(p7_mult_21_n880), .ZN(n853) );
  OAI21_X1 U1279 ( .B1(n852), .B2(p7_mult_21_n880), .A(p7_mult_21_n878), .ZN(
        n854) );
  AOI211_X1 U1280 ( .C1(n828), .C2(p7_mult_21_n889), .A(n873), .B(n851), .ZN(
        n852) );
  NAND2_X1 U1281 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U1282 ( .A1(p7_mult_21_n980), .A2(p7_mult_21_n981), .ZN(n858) );
  OAI21_X1 U1283 ( .B1(p7_mult_21_n980), .B2(p7_mult_21_n981), .A(
        p7_mult_21_n979), .ZN(n859) );
  NAND3_X1 U1284 ( .A1(n859), .A2(n858), .A3(p7_mult_21_n974), .ZN(n861) );
  AOI222_X1 U1285 ( .A1(p7_mult_21_n1040), .A2(p7_mult_21_n1041), .B1(n827), 
        .B2(p7_mult_21_n1040), .C1(n827), .C2(p7_mult_21_n1041), .ZN(
        p7_mult_21_n1034) );
  NAND2_X1 U1286 ( .A1(p7_mult_21_n1074), .A2(p7_mult_21_n1073), .ZN(n825) );
  NAND2_X1 U1287 ( .A1(p7_mult_21_n1074), .A2(p7_mult_21_n1075), .ZN(n823) );
  NAND2_X1 U1288 ( .A1(n844), .A2(p7_mult_21_n1149), .ZN(n868) );
  NAND2_X1 U1289 ( .A1(p7_mult_21_n1147), .A2(p7_mult_21_n1149), .ZN(n866) );
  NAND4_X1 U1290 ( .A1(n869), .A2(n868), .A3(p7_mult_21_n1108), .A4(n867), 
        .ZN(n871) );
  NAND4_X1 U1291 ( .A1(n866), .A2(n869), .A3(p7_mult_21_n1110), .A4(n867), 
        .ZN(n872) );
  NAND2_X1 U1292 ( .A1(n844), .A2(p7_mult_21_n1148), .ZN(n869) );
  AOI222_X1 U1293 ( .A1(p7_mult_21_n928), .A2(p7_mult_21_n929), .B1(
        p7_mult_21_n928), .B2(p7_mult_21_n930), .C1(p7_mult_21_n929), .C2(
        p7_mult_21_n930), .ZN(p7_mult_21_n895) );
  AOI221_X1 U1294 ( .B1(reg2_reg[9]), .B2(B1[0]), .C1(p7_mult_21_n945), .C2(
        n830), .A(p7_mult_21_n943), .ZN(p7_mult_21_n1333) );
  MUX2_X1 U1295 ( .A(p7_mult_21_n844), .B(p7_mult_21_n1262), .S(reg2_reg[0]), 
        .Z(p7_mult_21_n1247) );
  AOI221_X1 U1296 ( .B1(reg2_reg[11]), .B2(B1[0]), .C1(p7_mult_21_n911), .C2(
        n831), .A(p7_mult_21_n909), .ZN(p7_mult_21_n1398) );
  NAND2_X1 U1297 ( .A1(p7_mult_21_n1149), .A2(p7_mult_21_n1148), .ZN(n867) );
  NAND2_X1 U1298 ( .A1(p7_mult_21_n1108), .A2(p7_mult_21_n1110), .ZN(n870) );
  NAND2_X1 U1299 ( .A1(p7_mult_21_n972), .A2(p7_mult_21_n974), .ZN(n860) );
  XOR2_X1 U1300 ( .A(p7_mult_21_n900), .B(p7_mult_21_n913), .Z(p7_mult_21_n897) );
  AOI222_X1 U1301 ( .A1(p7_mult_21_n898), .A2(p7_mult_21_n899), .B1(
        p7_mult_21_n898), .B2(p7_mult_21_n900), .C1(p7_mult_21_n899), .C2(
        p7_mult_21_n900), .ZN(p7_mult_21_n889) );
  XOR2_X1 U1302 ( .A(p7_mult_21_n901), .B(p7_mult_21_n893), .Z(p7_mult_21_n891) );
  OAI21_X1 U1303 ( .B1(p7_mult_21_n867), .B2(p7_mult_21_n866), .A(
        p7_mult_21_n868), .ZN(n850) );
  AOI222_X1 U1304 ( .A1(p7_mult_21_n1147), .A2(p7_mult_21_n1148), .B1(
        p7_mult_21_n1147), .B2(p7_mult_21_n1149), .C1(p7_mult_21_n1148), .C2(
        p7_mult_21_n1149), .ZN(n843) );
  INV_X1 U1305 ( .A(p7_mult_21_n1095), .ZN(p7_mult_21_n1169) );
  INV_X1 U1306 ( .A(B1[3]), .ZN(n829) );
  INV_X1 U1307 ( .A(B1[2]), .ZN(n835) );
  INV_X1 U1308 ( .A(B1[1]), .ZN(n837) );
  INV_X1 U1309 ( .A(B1[1]), .ZN(n836) );
  INV_X1 U1310 ( .A(B1[2]), .ZN(p7_mult_21_n1180) );
  INV_X1 U1311 ( .A(B1[3]), .ZN(p7_mult_21_n1133) );
  INV_X1 U1312 ( .A(p7_mult_21_n1273), .ZN(p7_mult_21_n847) );
  INV_X1 U1313 ( .A(p7_mult_21_n1255), .ZN(p7_mult_21_n1254) );
  OR2_X1 U1314 ( .A1(p7_mult_21_n1253), .A2(p7_mult_21_n1252), .ZN(n822) );
  AND3_X1 U1315 ( .A1(n872), .A2(n871), .A3(n870), .ZN(p7_mult_21_n1074) );
  AND3_X1 U1316 ( .A1(n825), .A2(n823), .A3(n824), .ZN(n827) );
  AND2_X1 U1317 ( .A1(p7_mult_21_n980), .A2(p7_mult_21_n979), .ZN(n863) );
  AND2_X1 U1318 ( .A1(p7_mult_21_n980), .A2(p7_mult_21_n981), .ZN(n864) );
  AND2_X1 U1319 ( .A1(p7_mult_21_n979), .A2(p7_mult_21_n981), .ZN(n865) );
  AOI21_X1 U1320 ( .B1(n832), .B2(p7_mult_21_n972), .A(n862), .ZN(
        p7_mult_21_n933) );
  AND2_X1 U1321 ( .A1(p7_mult_21_n933), .A2(p7_mult_21_n934), .ZN(n855) );
  AND2_X1 U1322 ( .A1(p7_mult_21_n933), .A2(p7_mult_21_n932), .ZN(n856) );
  AND2_X1 U1323 ( .A1(p7_mult_21_n934), .A2(p7_mult_21_n932), .ZN(n857) );
  AND2_X1 U1324 ( .A1(p7_mult_21_n895), .A2(p7_mult_21_n896), .ZN(n840) );
  AND2_X1 U1325 ( .A1(p7_mult_21_n895), .A2(p7_mult_21_n897), .ZN(n839) );
  AND2_X1 U1326 ( .A1(p7_mult_21_n896), .A2(p7_mult_21_n897), .ZN(n838) );
  AND2_X1 U1327 ( .A1(p7_mult_21_n891), .A2(p7_mult_21_n889), .ZN(n873) );
  AND2_X1 U1328 ( .A1(p7_mult_21_n890), .A2(p7_mult_21_n891), .ZN(n851) );
  AND2_X1 U1329 ( .A1(n854), .A2(n853), .ZN(p7_mult_21_n865) );
  INV_X1 U1330 ( .A(p7_mult_21_n860), .ZN(n849) );
  NOR3_X2 U1331 ( .A1(n855), .A2(n856), .A3(n857), .ZN(p7_mult_21_n926) );
  AOI222_X4 U1332 ( .A1(p7_mult_21_n925), .A2(p7_mult_21_n926), .B1(
        p7_mult_21_n925), .B2(p7_mult_21_n927), .C1(p7_mult_21_n926), .C2(
        p7_mult_21_n927), .ZN(p7_mult_21_n896) );
  AOI222_X4 U1333 ( .A1(p7_mult_21_n1193), .A2(p7_mult_21_n1194), .B1(
        p7_mult_21_n1193), .B2(p7_mult_21_n1195), .C1(p7_mult_21_n1194), .C2(
        p7_mult_21_n1195), .ZN(p7_mult_21_n1183) );
  NOR3_X2 U1334 ( .A1(n840), .A2(n839), .A3(n838), .ZN(n828) );
  AOI221_X4 U1335 ( .B1(reg2_reg[2]), .B2(reg2_reg[3]), .C1(p7_mult_21_n1401), 
        .C2(p7_mult_21_n1126), .A(p7_mult_21_n1095), .ZN(p7_mult_21_n1096) );
  AND3_X2 U1336 ( .A1(n825), .A2(n823), .A3(n824), .ZN(p7_mult_21_n1042) );
  AOI222_X2 U1337 ( .A1(p7_mult_21_n1040), .A2(p7_mult_21_n1041), .B1(
        p7_mult_21_n1042), .B2(p7_mult_21_n1040), .C1(p7_mult_21_n1042), .C2(
        p7_mult_21_n1041), .ZN(n821) );
  AOI22_X1 U1338 ( .A1(reg2_reg[4]), .A2(reg2_reg[3]), .B1(p7_mult_21_n1126), 
        .B2(p7_mult_21_n1378), .ZN(p7_mult_21_n1028) );
  AOI221_X4 U1339 ( .B1(reg2_reg[4]), .B2(reg2_reg[5]), .C1(p7_mult_21_n1378), 
        .C2(p7_mult_21_n1053), .A(p7_mult_21_n1028), .ZN(p7_mult_21_n1029) );
  AOI222_X2 U1340 ( .A1(p7_mult_21_n1033), .A2(n821), .B1(p7_mult_21_n1033), 
        .B2(p7_mult_21_n1035), .C1(p7_mult_21_n1034), .C2(p7_mult_21_n1035), 
        .ZN(p7_mult_21_n980) );
  NOR3_X2 U1341 ( .A1(n863), .A2(n864), .A3(n865), .ZN(n832) );
  XNOR2_X1 U1342 ( .A(B0[2]), .B(reg1_reg[3]), .ZN(p6_mult_21_n709) );
  XNOR2_X1 U1343 ( .A(B0[1]), .B(reg1_reg[3]), .ZN(p6_mult_21_n708) );
  XNOR2_X1 U1344 ( .A(reg1_reg[3]), .B(B0[0]), .ZN(p6_mult_21_n705) );
  NOR2_X1 U1345 ( .A1(p6_mult_21_n722), .A2(p6_mult_21_n723), .ZN(
        p6_mult_21_n393) );
  XNOR2_X1 U1346 ( .A(B0[4]), .B(reg1_reg[3]), .ZN(p6_mult_21_n711) );
  XNOR2_X1 U1347 ( .A(B0[3]), .B(reg1_reg[3]), .ZN(p6_mult_21_n710) );
  OAI22_X1 U1348 ( .A1(p6_mult_21_n724), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n726), .ZN(p6_mult_21_n392) );
  XNOR2_X1 U1349 ( .A(B0[5]), .B(reg1_reg[3]), .ZN(p6_mult_21_n712) );
  OAI22_X1 U1350 ( .A1(p6_mult_21_n727), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n728), .ZN(p6_mult_21_n390) );
  XNOR2_X1 U1351 ( .A(B0[6]), .B(reg1_reg[3]), .ZN(p6_mult_21_n713) );
  OAI22_X1 U1352 ( .A1(p6_mult_21_n728), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n729), .ZN(p6_mult_21_n389) );
  XNOR2_X1 U1353 ( .A(B0[7]), .B(reg1_reg[3]), .ZN(p6_mult_21_n714) );
  XNOR2_X1 U1354 ( .A(B0[8]), .B(reg1_reg[3]), .ZN(p6_mult_21_n715) );
  OAI22_X1 U1355 ( .A1(p6_mult_21_n729), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n730), .ZN(p6_mult_21_n388) );
  XNOR2_X1 U1356 ( .A(B0[10]), .B(reg1_reg[3]), .ZN(p6_mult_21_n717) );
  XNOR2_X1 U1357 ( .A(B0[9]), .B(reg1_reg[3]), .ZN(p6_mult_21_n716) );
  OAI22_X1 U1358 ( .A1(p6_mult_21_n731), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n732), .ZN(p6_mult_21_n386) );
  OAI22_X1 U1359 ( .A1(p6_mult_21_n730), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n731), .ZN(p6_mult_21_n387) );
  XNOR2_X1 U1360 ( .A(B0[11]), .B(reg1_reg[3]), .ZN(p6_mult_21_n718) );
  OAI22_X1 U1361 ( .A1(p6_mult_21_n733), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n734), .ZN(p6_mult_21_n384) );
  XNOR2_X1 U1362 ( .A(B0[12]), .B(reg1_reg[3]), .ZN(p6_mult_21_n719) );
  OAI22_X1 U1363 ( .A1(p6_mult_21_n732), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n733), .ZN(p6_mult_21_n385) );
  XNOR2_X1 U1364 ( .A(B0[13]), .B(reg1_reg[3]), .ZN(p6_mult_21_n721) );
  NAND2_X1 U1365 ( .A1(p6_mult_21_n636), .A2(p6_mult_21_n299), .ZN(
        p6_mult_21_n642) );
  NAND2_X1 U1366 ( .A1(p6_mult_21_n636), .A2(p6_mult_21_n294), .ZN(
        p6_mult_21_n641) );
  OAI22_X1 U1367 ( .A1(p6_mult_21_n734), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n735), .ZN(p6_mult_21_n818) );
  OAI22_X1 U1368 ( .A1(p6_mult_21_n735), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n736), .ZN(p6_mult_21_n382) );
  OAI22_X1 U1369 ( .A1(p6_mult_21_n736), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n737), .ZN(p6_mult_21_n381) );
  NAND2_X1 U1370 ( .A1(p6_mult_21_n828), .A2(p6_mult_21_n277), .ZN(
        p6_mult_21_n679) );
  NAND2_X1 U1371 ( .A1(p6_mult_21_n828), .A2(p6_mult_21_n268), .ZN(
        p6_mult_21_n678) );
  OAI22_X1 U1372 ( .A1(p6_mult_21_n737), .A2(p6_mult_21_n725), .B1(
        p6_mult_21_n723), .B2(p6_mult_21_n739), .ZN(p6_mult_21_n209) );
  AOI21_X1 U1373 ( .B1(p6_mult_21_n725), .B2(p6_mult_21_n723), .A(
        p6_mult_21_n739), .ZN(p6_mult_21_n738) );
  OAI222_X1 U1374 ( .A1(p6_mult_21_n825), .A2(p6_mult_21_n826), .B1(
        p6_mult_21_n825), .B2(p6_mult_21_n827), .C1(p6_mult_21_n827), .C2(
        p6_mult_21_n826), .ZN(p6_mult_21_n640) );
  NAND2_X1 U1375 ( .A1(p6_mult_21_n640), .A2(p6_mult_21_n246), .ZN(
        p6_mult_21_n672) );
  NAND2_X1 U1376 ( .A1(n875), .A2(n874), .ZN(p6_mult_21_n140) );
  OAI21_X1 U1377 ( .B1(p6_mult_21_n174), .B2(p6_mult_21_n179), .A(
        p6_mult_21_n141), .ZN(n875) );
  NAND2_X1 U1378 ( .A1(n877), .A2(n876), .ZN(p6_mult_21_n141) );
  OAI21_X1 U1379 ( .B1(p6_mult_21_n185), .B2(p6_mult_21_n180), .A(
        p6_mult_21_n142), .ZN(n877) );
  NAND2_X1 U1380 ( .A1(n878), .A2(p6_mult_21_n234), .ZN(n879) );
  NAND2_X1 U1381 ( .A1(p6_mult_21_n148), .A2(p6_mult_21_n245), .ZN(n881) );
  NAND3_X1 U1382 ( .A1(p6_mult_21_n672), .A2(p6_mult_21_n673), .A3(
        p6_mult_21_n674), .ZN(n878) );
  NAND3_X1 U1383 ( .A1(n881), .A2(n880), .A3(n879), .ZN(p6_mult_21_n147) );
  NAND2_X1 U1384 ( .A1(p6_mult_21_n234), .A2(p6_mult_21_n245), .ZN(n880) );
  NAND2_X1 U1385 ( .A1(p6_mult_21_n180), .A2(p6_mult_21_n185), .ZN(n876) );
  NAND2_X1 U1386 ( .A1(p6_mult_21_n174), .A2(p6_mult_21_n179), .ZN(n874) );
  OR3_X1 U1387 ( .A1(p6_mult_21_n723), .A2(B0[0]), .A3(p6_mult_21_n807), .ZN(
        p6_mult_21_n808) );
  INV_X1 U1388 ( .A(VIN), .ZN(n940) );
  INV_X1 U1389 ( .A(VIN), .ZN(n941) );
  OR2_X1 U1390 ( .A1(VIN), .A2(SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_), 
        .ZN(n935) );
  OR2_X1 U1391 ( .A1(VIN), .A2(n918), .ZN(n934) );
  INV_X1 U1392 ( .A(VIN), .ZN(n942) );
  NAND2_X1 U1393 ( .A1(temp5[11]), .A2(VIN), .ZN(n936) );
  NAND2_X1 U1394 ( .A1(n936), .A2(n935), .ZN(REG51_n255) );
  NAND2_X1 U1395 ( .A1(temp2[13]), .A2(VIN), .ZN(REG2_1_n75) );
  NAND2_X1 U1396 ( .A1(temp4[12]), .A2(VIN), .ZN(n937) );
  NAND2_X1 U1397 ( .A1(n937), .A2(n934), .ZN(REG4_1_n254) );
  MUX2_X1 U1398 ( .A(temp4[13]), .B(mul4_reg[13]), .S(n942), .Z(REG4_1_n253)
         );
  NAND2_X1 U1399 ( .A1(reg6[13]), .A2(n942), .ZN(n939) );
  NAND2_X1 U1400 ( .A1(temp5[13]), .A2(VIN), .ZN(n938) );
  NAND2_X1 U1401 ( .A1(n938), .A2(n939), .ZN(REG51_n253) );
  OAI21_X1 U1402 ( .B1(VIN), .B2(n889), .A(n286), .ZN(REG31_n263) );
  NAND2_X1 U1403 ( .A1(n286), .A2(n287), .ZN(REGISTER2_n263) );
  OAI22_X1 U1404 ( .A1(n941), .A2(reg4[1]), .B1(reg5[1]), .B2(VIN), .ZN(n315)
         );
endmodule

