
module IIR_CA ( CLK, RST_n, VIN, DIN, B0, B1, B2, A1, A2, VOUT, DOUT );
  input [13:0] DIN;
  input [13:0] B0;
  input [13:0] B1;
  input [13:0] B2;
  input [13:0] A1;
  input [13:0] A2;
  output [13:0] DOUT;
  input CLK, RST_n, VIN;
  output VOUT;
  wire   n2, n3, n6, n7, n10, n11, n14, n15, n18, n19, n22, n23, n26, n27, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, temp5_26_,
         temp5_25_, temp5_24_, temp5_23_, temp5_22_, temp5_21_, temp5_20_,
         temp5_19_, temp5_18_, temp5_17_, temp5_16_, temp5_15_, temp5_14_,
         temp5_13_, temp4_26_, temp4_25_, temp4_24_, temp4_23_, temp4_22_,
         temp4_21_, temp4_20_, temp4_19_, temp4_18_, temp4_17_, temp4_16_,
         temp4_15_, temp4_14_, temp4_13_, temp3_26_, temp3_25_, temp3_24_,
         temp3_23_, temp3_22_, temp3_21_, temp3_20_, temp3_19_, temp3_18_,
         temp3_17_, temp3_16_, temp3_15_, temp3_14_, temp3_13_, ff_9_, ff_8_,
         ff_7_, ff_6_, ff_5_, ff_4_, ff_3_, ff_2_, ff_1_, ff_13_, ff_12_,
         ff_11_, ff_10_, ff_0_, temp2_26_, temp2_25_, temp2_24_, temp2_23_,
         temp2_22_, temp2_21_, temp2_20_, temp2_19_, temp2_18_, temp2_17_,
         temp2_16_, temp2_15_, temp2_14_, temp2_13_, temp1_26_, temp1_25_,
         temp1_24_, temp1_23_, temp1_22_, temp1_21_, temp1_20_, temp1_19_,
         temp1_18_, temp1_17_, temp1_16_, temp1_15_, temp1_14_, temp1_13_,
         fb_9_, fb_8_, fb_7_, fb_6_, fb_5_, fb_4_, fb_3_, fb_2_, fb_1_, fb_13_,
         fb_12_, fb_11_, fb_10_, fb_0_, N9, N8, N7, N6, N5, N4, N3, N2, N13,
         N12, N11, N10, N1, N0, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, mult_50_n805, mult_50_n804,
         mult_50_n803, mult_50_n802, mult_50_n801, mult_50_n800, mult_50_n799,
         mult_50_n798, mult_50_n797, mult_50_n796, mult_50_n795, mult_50_n794,
         mult_50_n793, mult_50_n792, mult_50_n791, mult_50_n790, mult_50_n789,
         mult_50_n788, mult_50_n787, mult_50_n786, mult_50_n785, mult_50_n784,
         mult_50_n783, mult_50_n782, mult_50_n781, mult_50_n780, mult_50_n779,
         mult_50_n778, mult_50_n777, mult_50_n776, mult_50_n775, mult_50_n774,
         mult_50_n773, mult_50_n772, mult_50_n771, mult_50_n770, mult_50_n769,
         mult_50_n768, mult_50_n767, mult_50_n766, mult_50_n765, mult_50_n764,
         mult_50_n763, mult_50_n762, mult_50_n761, mult_50_n760, mult_50_n759,
         mult_50_n758, mult_50_n757, mult_50_n756, mult_50_n755, mult_50_n754,
         mult_50_n753, mult_50_n752, mult_50_n751, mult_50_n750, mult_50_n749,
         mult_50_n748, mult_50_n747, mult_50_n746, mult_50_n745, mult_50_n744,
         mult_50_n743, mult_50_n742, mult_50_n741, mult_50_n740, mult_50_n739,
         mult_50_n738, mult_50_n737, mult_50_n736, mult_50_n735, mult_50_n734,
         mult_50_n733, mult_50_n732, mult_50_n731, mult_50_n730, mult_50_n729,
         mult_50_n728, mult_50_n727, mult_50_n726, mult_50_n725, mult_50_n724,
         mult_50_n723, mult_50_n722, mult_50_n721, mult_50_n720, mult_50_n719,
         mult_50_n718, mult_50_n717, mult_50_n716, mult_50_n715, mult_50_n714,
         mult_50_n713, mult_50_n712, mult_50_n711, mult_50_n710, mult_50_n709,
         mult_50_n708, mult_50_n707, mult_50_n706, mult_50_n705, mult_50_n704,
         mult_50_n703, mult_50_n702, mult_50_n701, mult_50_n700, mult_50_n699,
         mult_50_n698, mult_50_n697, mult_50_n696, mult_50_n695, mult_50_n694,
         mult_50_n693, mult_50_n692, mult_50_n691, mult_50_n690, mult_50_n689,
         mult_50_n688, mult_50_n687, mult_50_n686, mult_50_n685, mult_50_n684,
         mult_50_n683, mult_50_n682, mult_50_n681, mult_50_n680, mult_50_n679,
         mult_50_n678, mult_50_n677, mult_50_n676, mult_50_n675, mult_50_n674,
         mult_50_n673, mult_50_n672, mult_50_n671, mult_50_n670, mult_50_n669,
         mult_50_n668, mult_50_n667, mult_50_n666, mult_50_n665, mult_50_n664,
         mult_50_n663, mult_50_n662, mult_50_n661, mult_50_n660, mult_50_n659,
         mult_50_n658, mult_50_n657, mult_50_n656, mult_50_n655, mult_50_n654,
         mult_50_n653, mult_50_n652, mult_50_n651, mult_50_n650, mult_50_n649,
         mult_50_n648, mult_50_n647, mult_50_n646, mult_50_n645, mult_50_n644,
         mult_50_n643, mult_50_n642, mult_50_n641, mult_50_n640, mult_50_n639,
         mult_50_n638, mult_50_n637, mult_50_n636, mult_50_n635, mult_50_n419,
         mult_50_n418, mult_50_n417, mult_50_n416, mult_50_n415, mult_50_n414,
         mult_50_n413, mult_50_n412, mult_50_n411, mult_50_n410, mult_50_n409,
         mult_50_n408, mult_50_n406, mult_50_n405, mult_50_n404, mult_50_n403,
         mult_50_n402, mult_50_n401, mult_50_n400, mult_50_n399, mult_50_n398,
         mult_50_n397, mult_50_n396, mult_50_n395, mult_50_n394, mult_50_n393,
         mult_50_n392, mult_50_n391, mult_50_n390, mult_50_n389, mult_50_n388,
         mult_50_n387, mult_50_n386, mult_50_n385, mult_50_n384, mult_50_n382,
         mult_50_n381, mult_50_n380, mult_50_n379, mult_50_n378, mult_50_n377,
         mult_50_n376, mult_50_n375, mult_50_n374, mult_50_n373, mult_50_n372,
         mult_50_n371, mult_50_n370, mult_50_n369, mult_50_n368, mult_50_n367,
         mult_50_n366, mult_50_n365, mult_50_n364, mult_50_n363, mult_50_n362,
         mult_50_n361, mult_50_n360, mult_50_n359, mult_50_n358, mult_50_n357,
         mult_50_n356, mult_50_n355, mult_50_n354, mult_50_n353, mult_50_n352,
         mult_50_n351, mult_50_n350, mult_50_n349, mult_50_n348, mult_50_n346,
         mult_50_n345, mult_50_n344, mult_50_n343, mult_50_n342, mult_50_n341,
         mult_50_n340, mult_50_n339, mult_50_n338, mult_50_n337, mult_50_n336,
         mult_50_n335, mult_50_n334, mult_50_n333, mult_50_n332, mult_50_n331,
         mult_50_n330, mult_50_n329, mult_50_n328, mult_50_n327, mult_50_n326,
         mult_50_n325, mult_50_n321, mult_50_n320, mult_50_n319, mult_50_n318,
         mult_50_n317, mult_50_n316, mult_50_n315, mult_50_n314, mult_50_n313,
         mult_50_n312, mult_50_n311, mult_50_n310, mult_50_n309, mult_50_n308,
         mult_50_n307, mult_50_n306, mult_50_n305, mult_50_n304, mult_50_n303,
         mult_50_n302, mult_50_n301, mult_50_n300, mult_50_n299, mult_50_n298,
         mult_50_n297, mult_50_n296, mult_50_n295, mult_50_n294, mult_50_n293,
         mult_50_n292, mult_50_n291, mult_50_n290, mult_50_n289, mult_50_n288,
         mult_50_n287, mult_50_n286, mult_50_n285, mult_50_n284, mult_50_n283,
         mult_50_n282, mult_50_n281, mult_50_n280, mult_50_n279, mult_50_n278,
         mult_50_n277, mult_50_n276, mult_50_n275, mult_50_n274, mult_50_n273,
         mult_50_n272, mult_50_n271, mult_50_n270, mult_50_n269, mult_50_n268,
         mult_50_n267, mult_50_n266, mult_50_n265, mult_50_n264, mult_50_n263,
         mult_50_n262, mult_50_n261, mult_50_n260, mult_50_n259, mult_50_n258,
         mult_50_n257, mult_50_n256, mult_50_n255, mult_50_n254, mult_50_n253,
         mult_50_n252, mult_50_n251, mult_50_n250, mult_50_n249, mult_50_n248,
         mult_50_n247, mult_50_n246, mult_50_n245, mult_50_n244, mult_50_n243,
         mult_50_n242, mult_50_n241, mult_50_n240, mult_50_n239, mult_50_n238,
         mult_50_n237, mult_50_n236, mult_50_n235, mult_50_n234, mult_50_n233,
         mult_50_n232, mult_50_n231, mult_50_n230, mult_50_n229, mult_50_n228,
         mult_50_n227, mult_50_n226, mult_50_n225, mult_50_n224, mult_50_n223,
         mult_50_n222, mult_50_n221, mult_50_n220, mult_50_n219, mult_50_n218,
         mult_50_n217, mult_50_n216, mult_50_n215, mult_50_n214, mult_50_n213,
         mult_50_n212, mult_50_n211, mult_50_n210, mult_50_n209, mult_50_n208,
         mult_50_n207, mult_50_n206, mult_50_n205, mult_50_n204, mult_50_n203,
         mult_50_n202, mult_50_n201, mult_50_n200, mult_50_n199, mult_50_n198,
         mult_50_n197, mult_50_n196, mult_50_n195, mult_50_n194, mult_50_n193,
         mult_50_n192, mult_50_n191, mult_50_n190, mult_50_n189, mult_50_n188,
         mult_50_n187, mult_50_n186, mult_50_n185, mult_50_n184, mult_50_n183,
         mult_50_n182, mult_50_n181, mult_50_n180, mult_50_n179, mult_50_n178,
         mult_50_n177, mult_50_n176, mult_50_n175, mult_50_n174, mult_50_n173,
         mult_50_n172, mult_50_n171, mult_50_n170, mult_50_n169, mult_50_n168,
         mult_50_n167, mult_50_n166, mult_50_n165, mult_50_n164, mult_50_n163,
         mult_50_n162, mult_50_n149, mult_50_n148, mult_50_n147, mult_50_n146,
         mult_50_n145, mult_50_n144, mult_50_n143, mult_50_n142, mult_50_n141,
         mult_50_n140, mult_50_n139, mult_50_n138, mult_50_n137, mult_50_n136,
         mult_52_n805, mult_52_n804, mult_52_n803, mult_52_n802, mult_52_n801,
         mult_52_n800, mult_52_n799, mult_52_n798, mult_52_n797, mult_52_n796,
         mult_52_n795, mult_52_n794, mult_52_n793, mult_52_n792, mult_52_n791,
         mult_52_n790, mult_52_n789, mult_52_n788, mult_52_n787, mult_52_n786,
         mult_52_n785, mult_52_n784, mult_52_n783, mult_52_n782, mult_52_n781,
         mult_52_n780, mult_52_n779, mult_52_n778, mult_52_n777, mult_52_n776,
         mult_52_n775, mult_52_n774, mult_52_n773, mult_52_n772, mult_52_n771,
         mult_52_n770, mult_52_n769, mult_52_n768, mult_52_n767, mult_52_n766,
         mult_52_n765, mult_52_n764, mult_52_n763, mult_52_n762, mult_52_n761,
         mult_52_n760, mult_52_n759, mult_52_n758, mult_52_n757, mult_52_n756,
         mult_52_n755, mult_52_n754, mult_52_n753, mult_52_n752, mult_52_n751,
         mult_52_n750, mult_52_n749, mult_52_n748, mult_52_n747, mult_52_n746,
         mult_52_n745, mult_52_n744, mult_52_n743, mult_52_n742, mult_52_n741,
         mult_52_n740, mult_52_n739, mult_52_n738, mult_52_n737, mult_52_n736,
         mult_52_n735, mult_52_n734, mult_52_n733, mult_52_n732, mult_52_n731,
         mult_52_n730, mult_52_n729, mult_52_n728, mult_52_n727, mult_52_n726,
         mult_52_n725, mult_52_n724, mult_52_n723, mult_52_n722, mult_52_n721,
         mult_52_n720, mult_52_n719, mult_52_n718, mult_52_n717, mult_52_n716,
         mult_52_n715, mult_52_n714, mult_52_n713, mult_52_n712, mult_52_n711,
         mult_52_n710, mult_52_n709, mult_52_n708, mult_52_n707, mult_52_n706,
         mult_52_n705, mult_52_n704, mult_52_n703, mult_52_n702, mult_52_n701,
         mult_52_n700, mult_52_n699, mult_52_n698, mult_52_n697, mult_52_n696,
         mult_52_n695, mult_52_n694, mult_52_n693, mult_52_n692, mult_52_n691,
         mult_52_n690, mult_52_n689, mult_52_n688, mult_52_n687, mult_52_n686,
         mult_52_n685, mult_52_n684, mult_52_n683, mult_52_n682, mult_52_n681,
         mult_52_n680, mult_52_n679, mult_52_n678, mult_52_n677, mult_52_n676,
         mult_52_n675, mult_52_n674, mult_52_n673, mult_52_n672, mult_52_n671,
         mult_52_n670, mult_52_n669, mult_52_n668, mult_52_n667, mult_52_n666,
         mult_52_n665, mult_52_n664, mult_52_n663, mult_52_n662, mult_52_n661,
         mult_52_n660, mult_52_n659, mult_52_n658, mult_52_n657, mult_52_n656,
         mult_52_n655, mult_52_n654, mult_52_n653, mult_52_n652, mult_52_n651,
         mult_52_n650, mult_52_n649, mult_52_n648, mult_52_n647, mult_52_n646,
         mult_52_n645, mult_52_n644, mult_52_n643, mult_52_n642, mult_52_n641,
         mult_52_n640, mult_52_n639, mult_52_n638, mult_52_n637, mult_52_n636,
         mult_52_n635, mult_52_n419, mult_52_n418, mult_52_n417, mult_52_n416,
         mult_52_n415, mult_52_n414, mult_52_n413, mult_52_n412, mult_52_n411,
         mult_52_n410, mult_52_n409, mult_52_n408, mult_52_n406, mult_52_n405,
         mult_52_n404, mult_52_n403, mult_52_n402, mult_52_n401, mult_52_n400,
         mult_52_n399, mult_52_n398, mult_52_n397, mult_52_n396, mult_52_n395,
         mult_52_n394, mult_52_n393, mult_52_n392, mult_52_n391, mult_52_n390,
         mult_52_n389, mult_52_n388, mult_52_n387, mult_52_n386, mult_52_n385,
         mult_52_n384, mult_52_n382, mult_52_n381, mult_52_n380, mult_52_n379,
         mult_52_n378, mult_52_n377, mult_52_n376, mult_52_n375, mult_52_n374,
         mult_52_n373, mult_52_n372, mult_52_n371, mult_52_n370, mult_52_n369,
         mult_52_n368, mult_52_n367, mult_52_n366, mult_52_n365, mult_52_n364,
         mult_52_n363, mult_52_n362, mult_52_n361, mult_52_n360, mult_52_n359,
         mult_52_n358, mult_52_n357, mult_52_n356, mult_52_n355, mult_52_n354,
         mult_52_n353, mult_52_n352, mult_52_n351, mult_52_n350, mult_52_n349,
         mult_52_n348, mult_52_n346, mult_52_n345, mult_52_n344, mult_52_n343,
         mult_52_n342, mult_52_n341, mult_52_n340, mult_52_n339, mult_52_n338,
         mult_52_n337, mult_52_n336, mult_52_n335, mult_52_n334, mult_52_n333,
         mult_52_n332, mult_52_n331, mult_52_n330, mult_52_n329, mult_52_n328,
         mult_52_n327, mult_52_n326, mult_52_n325, mult_52_n321, mult_52_n320,
         mult_52_n319, mult_52_n318, mult_52_n317, mult_52_n316, mult_52_n315,
         mult_52_n314, mult_52_n313, mult_52_n312, mult_52_n311, mult_52_n310,
         mult_52_n309, mult_52_n308, mult_52_n307, mult_52_n306, mult_52_n305,
         mult_52_n304, mult_52_n303, mult_52_n302, mult_52_n301, mult_52_n300,
         mult_52_n299, mult_52_n298, mult_52_n297, mult_52_n296, mult_52_n295,
         mult_52_n294, mult_52_n293, mult_52_n292, mult_52_n291, mult_52_n290,
         mult_52_n289, mult_52_n288, mult_52_n287, mult_52_n286, mult_52_n285,
         mult_52_n284, mult_52_n283, mult_52_n282, mult_52_n281, mult_52_n280,
         mult_52_n279, mult_52_n278, mult_52_n277, mult_52_n276, mult_52_n275,
         mult_52_n274, mult_52_n273, mult_52_n272, mult_52_n271, mult_52_n270,
         mult_52_n269, mult_52_n268, mult_52_n267, mult_52_n266, mult_52_n265,
         mult_52_n264, mult_52_n263, mult_52_n262, mult_52_n261, mult_52_n260,
         mult_52_n259, mult_52_n258, mult_52_n257, mult_52_n256, mult_52_n255,
         mult_52_n254, mult_52_n253, mult_52_n252, mult_52_n251, mult_52_n250,
         mult_52_n249, mult_52_n248, mult_52_n247, mult_52_n246, mult_52_n245,
         mult_52_n244, mult_52_n243, mult_52_n242, mult_52_n241, mult_52_n240,
         mult_52_n239, mult_52_n238, mult_52_n237, mult_52_n236, mult_52_n235,
         mult_52_n234, mult_52_n233, mult_52_n232, mult_52_n231, mult_52_n230,
         mult_52_n229, mult_52_n228, mult_52_n227, mult_52_n226, mult_52_n225,
         mult_52_n224, mult_52_n223, mult_52_n222, mult_52_n221, mult_52_n220,
         mult_52_n219, mult_52_n218, mult_52_n217, mult_52_n216, mult_52_n215,
         mult_52_n214, mult_52_n213, mult_52_n212, mult_52_n211, mult_52_n210,
         mult_52_n209, mult_52_n208, mult_52_n207, mult_52_n206, mult_52_n205,
         mult_52_n204, mult_52_n203, mult_52_n202, mult_52_n201, mult_52_n200,
         mult_52_n199, mult_52_n198, mult_52_n197, mult_52_n196, mult_52_n195,
         mult_52_n194, mult_52_n193, mult_52_n192, mult_52_n191, mult_52_n190,
         mult_52_n189, mult_52_n188, mult_52_n187, mult_52_n186, mult_52_n185,
         mult_52_n184, mult_52_n183, mult_52_n182, mult_52_n181, mult_52_n180,
         mult_52_n179, mult_52_n178, mult_52_n177, mult_52_n176, mult_52_n175,
         mult_52_n174, mult_52_n173, mult_52_n172, mult_52_n171, mult_52_n170,
         mult_52_n169, mult_52_n168, mult_52_n167, mult_52_n166, mult_52_n165,
         mult_52_n164, mult_52_n163, mult_52_n162, mult_52_n149, mult_52_n148,
         mult_52_n147, mult_52_n146, mult_52_n145, mult_52_n144, mult_52_n143,
         mult_52_n142, mult_52_n141, mult_52_n140, mult_52_n139, mult_52_n138,
         mult_52_n137, mult_52_n136, add_1_root_add_0_root_add_59_carry_1_,
         add_1_root_add_0_root_add_59_carry_2_,
         add_1_root_add_0_root_add_59_carry_3_,
         add_1_root_add_0_root_add_59_carry_4_,
         add_1_root_add_0_root_add_59_carry_5_,
         add_1_root_add_0_root_add_59_carry_6_,
         add_1_root_add_0_root_add_59_carry_7_,
         add_1_root_add_0_root_add_59_carry_8_,
         add_1_root_add_0_root_add_59_carry_9_,
         add_1_root_add_0_root_add_59_carry_10_,
         add_1_root_add_0_root_add_59_carry_11_,
         add_1_root_add_0_root_add_59_carry_12_,
         add_1_root_add_0_root_add_59_carry_13_, mult_54_n805, mult_54_n804,
         mult_54_n803, mult_54_n802, mult_54_n801, mult_54_n800, mult_54_n799,
         mult_54_n798, mult_54_n797, mult_54_n796, mult_54_n795, mult_54_n794,
         mult_54_n793, mult_54_n792, mult_54_n791, mult_54_n790, mult_54_n789,
         mult_54_n788, mult_54_n787, mult_54_n786, mult_54_n785, mult_54_n784,
         mult_54_n783, mult_54_n782, mult_54_n781, mult_54_n780, mult_54_n779,
         mult_54_n778, mult_54_n777, mult_54_n776, mult_54_n775, mult_54_n774,
         mult_54_n773, mult_54_n772, mult_54_n771, mult_54_n770, mult_54_n769,
         mult_54_n768, mult_54_n767, mult_54_n766, mult_54_n765, mult_54_n764,
         mult_54_n763, mult_54_n762, mult_54_n761, mult_54_n760, mult_54_n759,
         mult_54_n758, mult_54_n757, mult_54_n756, mult_54_n755, mult_54_n754,
         mult_54_n753, mult_54_n752, mult_54_n751, mult_54_n750, mult_54_n749,
         mult_54_n748, mult_54_n747, mult_54_n746, mult_54_n745, mult_54_n744,
         mult_54_n743, mult_54_n742, mult_54_n741, mult_54_n740, mult_54_n739,
         mult_54_n738, mult_54_n737, mult_54_n736, mult_54_n735, mult_54_n734,
         mult_54_n733, mult_54_n732, mult_54_n731, mult_54_n730, mult_54_n729,
         mult_54_n728, mult_54_n727, mult_54_n726, mult_54_n725, mult_54_n724,
         mult_54_n723, mult_54_n722, mult_54_n721, mult_54_n720, mult_54_n719,
         mult_54_n718, mult_54_n717, mult_54_n716, mult_54_n715, mult_54_n714,
         mult_54_n713, mult_54_n712, mult_54_n711, mult_54_n710, mult_54_n709,
         mult_54_n708, mult_54_n707, mult_54_n706, mult_54_n705, mult_54_n704,
         mult_54_n703, mult_54_n702, mult_54_n701, mult_54_n700, mult_54_n699,
         mult_54_n698, mult_54_n697, mult_54_n696, mult_54_n695, mult_54_n694,
         mult_54_n693, mult_54_n692, mult_54_n691, mult_54_n690, mult_54_n689,
         mult_54_n688, mult_54_n687, mult_54_n686, mult_54_n685, mult_54_n684,
         mult_54_n683, mult_54_n682, mult_54_n681, mult_54_n680, mult_54_n679,
         mult_54_n678, mult_54_n677, mult_54_n676, mult_54_n675, mult_54_n674,
         mult_54_n673, mult_54_n672, mult_54_n671, mult_54_n670, mult_54_n669,
         mult_54_n668, mult_54_n667, mult_54_n666, mult_54_n665, mult_54_n664,
         mult_54_n663, mult_54_n662, mult_54_n661, mult_54_n660, mult_54_n659,
         mult_54_n658, mult_54_n657, mult_54_n656, mult_54_n655, mult_54_n654,
         mult_54_n653, mult_54_n652, mult_54_n651, mult_54_n650, mult_54_n649,
         mult_54_n648, mult_54_n647, mult_54_n646, mult_54_n645, mult_54_n644,
         mult_54_n643, mult_54_n642, mult_54_n641, mult_54_n640, mult_54_n639,
         mult_54_n638, mult_54_n637, mult_54_n636, mult_54_n635, mult_54_n419,
         mult_54_n418, mult_54_n417, mult_54_n416, mult_54_n415, mult_54_n414,
         mult_54_n413, mult_54_n412, mult_54_n411, mult_54_n410, mult_54_n409,
         mult_54_n408, mult_54_n406, mult_54_n405, mult_54_n404, mult_54_n403,
         mult_54_n402, mult_54_n401, mult_54_n400, mult_54_n399, mult_54_n398,
         mult_54_n397, mult_54_n396, mult_54_n395, mult_54_n394, mult_54_n393,
         mult_54_n392, mult_54_n391, mult_54_n390, mult_54_n389, mult_54_n388,
         mult_54_n387, mult_54_n386, mult_54_n385, mult_54_n384, mult_54_n382,
         mult_54_n381, mult_54_n380, mult_54_n379, mult_54_n378, mult_54_n377,
         mult_54_n376, mult_54_n375, mult_54_n374, mult_54_n373, mult_54_n372,
         mult_54_n371, mult_54_n370, mult_54_n369, mult_54_n368, mult_54_n367,
         mult_54_n366, mult_54_n365, mult_54_n364, mult_54_n363, mult_54_n362,
         mult_54_n361, mult_54_n360, mult_54_n359, mult_54_n358, mult_54_n357,
         mult_54_n356, mult_54_n355, mult_54_n354, mult_54_n353, mult_54_n352,
         mult_54_n351, mult_54_n350, mult_54_n349, mult_54_n348, mult_54_n346,
         mult_54_n345, mult_54_n344, mult_54_n343, mult_54_n342, mult_54_n341,
         mult_54_n340, mult_54_n339, mult_54_n338, mult_54_n337, mult_54_n336,
         mult_54_n335, mult_54_n334, mult_54_n333, mult_54_n332, mult_54_n331,
         mult_54_n330, mult_54_n329, mult_54_n328, mult_54_n327, mult_54_n326,
         mult_54_n325, mult_54_n321, mult_54_n320, mult_54_n319, mult_54_n318,
         mult_54_n317, mult_54_n316, mult_54_n315, mult_54_n314, mult_54_n313,
         mult_54_n312, mult_54_n311, mult_54_n310, mult_54_n309, mult_54_n308,
         mult_54_n307, mult_54_n306, mult_54_n305, mult_54_n304, mult_54_n303,
         mult_54_n302, mult_54_n301, mult_54_n300, mult_54_n299, mult_54_n298,
         mult_54_n297, mult_54_n296, mult_54_n295, mult_54_n294, mult_54_n293,
         mult_54_n292, mult_54_n291, mult_54_n290, mult_54_n289, mult_54_n288,
         mult_54_n287, mult_54_n286, mult_54_n285, mult_54_n284, mult_54_n283,
         mult_54_n282, mult_54_n281, mult_54_n280, mult_54_n279, mult_54_n278,
         mult_54_n277, mult_54_n276, mult_54_n275, mult_54_n274, mult_54_n273,
         mult_54_n272, mult_54_n271, mult_54_n270, mult_54_n269, mult_54_n268,
         mult_54_n267, mult_54_n266, mult_54_n265, mult_54_n264, mult_54_n263,
         mult_54_n262, mult_54_n261, mult_54_n260, mult_54_n259, mult_54_n258,
         mult_54_n257, mult_54_n256, mult_54_n255, mult_54_n254, mult_54_n253,
         mult_54_n252, mult_54_n251, mult_54_n250, mult_54_n249, mult_54_n248,
         mult_54_n247, mult_54_n246, mult_54_n245, mult_54_n244, mult_54_n243,
         mult_54_n242, mult_54_n241, mult_54_n240, mult_54_n239, mult_54_n238,
         mult_54_n237, mult_54_n236, mult_54_n235, mult_54_n234, mult_54_n233,
         mult_54_n232, mult_54_n231, mult_54_n230, mult_54_n229, mult_54_n228,
         mult_54_n227, mult_54_n226, mult_54_n225, mult_54_n224, mult_54_n223,
         mult_54_n222, mult_54_n221, mult_54_n220, mult_54_n219, mult_54_n218,
         mult_54_n217, mult_54_n216, mult_54_n215, mult_54_n214, mult_54_n213,
         mult_54_n212, mult_54_n211, mult_54_n210, mult_54_n209, mult_54_n208,
         mult_54_n207, mult_54_n206, mult_54_n205, mult_54_n204, mult_54_n203,
         mult_54_n202, mult_54_n201, mult_54_n200, mult_54_n199, mult_54_n198,
         mult_54_n197, mult_54_n196, mult_54_n195, mult_54_n194, mult_54_n193,
         mult_54_n192, mult_54_n191, mult_54_n190, mult_54_n189, mult_54_n188,
         mult_54_n187, mult_54_n186, mult_54_n185, mult_54_n184, mult_54_n183,
         mult_54_n182, mult_54_n181, mult_54_n180, mult_54_n179, mult_54_n178,
         mult_54_n177, mult_54_n176, mult_54_n175, mult_54_n174, mult_54_n173,
         mult_54_n172, mult_54_n171, mult_54_n170, mult_54_n169, mult_54_n168,
         mult_54_n167, mult_54_n166, mult_54_n165, mult_54_n164, mult_54_n163,
         mult_54_n162, mult_54_n149, mult_54_n148, mult_54_n147, mult_54_n146,
         mult_54_n145, mult_54_n144, mult_54_n143, mult_54_n142, mult_54_n141,
         mult_54_n140, mult_54_n139, mult_54_n138, mult_54_n137, mult_54_n136,
         add_0_root_add_0_root_add_59_carry_1_,
         add_0_root_add_0_root_add_59_carry_2_,
         add_0_root_add_0_root_add_59_carry_3_,
         add_0_root_add_0_root_add_59_carry_4_,
         add_0_root_add_0_root_add_59_carry_5_,
         add_0_root_add_0_root_add_59_carry_6_,
         add_0_root_add_0_root_add_59_carry_7_,
         add_0_root_add_0_root_add_59_carry_8_,
         add_0_root_add_0_root_add_59_carry_9_,
         add_0_root_add_0_root_add_59_carry_10_,
         add_0_root_add_0_root_add_59_carry_11_,
         add_0_root_add_0_root_add_59_carry_12_,
         add_0_root_add_0_root_add_59_carry_13_, mult_46_n812, mult_46_n811,
         mult_46_n810, mult_46_n809, mult_46_n808, mult_46_n807, mult_46_n806,
         mult_46_n805, mult_46_n804, mult_46_n803, mult_46_n802, mult_46_n801,
         mult_46_n800, mult_46_n799, mult_46_n798, mult_46_n797, mult_46_n796,
         mult_46_n795, mult_46_n794, mult_46_n793, mult_46_n792, mult_46_n791,
         mult_46_n790, mult_46_n789, mult_46_n788, mult_46_n787, mult_46_n786,
         mult_46_n785, mult_46_n784, mult_46_n783, mult_46_n782, mult_46_n781,
         mult_46_n780, mult_46_n779, mult_46_n778, mult_46_n777, mult_46_n776,
         mult_46_n775, mult_46_n774, mult_46_n773, mult_46_n772, mult_46_n771,
         mult_46_n770, mult_46_n769, mult_46_n768, mult_46_n767, mult_46_n766,
         mult_46_n765, mult_46_n764, mult_46_n763, mult_46_n762, mult_46_n761,
         mult_46_n760, mult_46_n759, mult_46_n758, mult_46_n757, mult_46_n756,
         mult_46_n755, mult_46_n754, mult_46_n753, mult_46_n752, mult_46_n751,
         mult_46_n750, mult_46_n749, mult_46_n748, mult_46_n747, mult_46_n746,
         mult_46_n745, mult_46_n744, mult_46_n743, mult_46_n742, mult_46_n741,
         mult_46_n740, mult_46_n739, mult_46_n738, mult_46_n737, mult_46_n736,
         mult_46_n735, mult_46_n734, mult_46_n733, mult_46_n732, mult_46_n731,
         mult_46_n730, mult_46_n729, mult_46_n728, mult_46_n727, mult_46_n726,
         mult_46_n725, mult_46_n724, mult_46_n723, mult_46_n722, mult_46_n721,
         mult_46_n720, mult_46_n719, mult_46_n718, mult_46_n717, mult_46_n716,
         mult_46_n715, mult_46_n714, mult_46_n713, mult_46_n712, mult_46_n711,
         mult_46_n710, mult_46_n709, mult_46_n708, mult_46_n707, mult_46_n706,
         mult_46_n705, mult_46_n704, mult_46_n703, mult_46_n702, mult_46_n701,
         mult_46_n700, mult_46_n699, mult_46_n698, mult_46_n697, mult_46_n696,
         mult_46_n695, mult_46_n694, mult_46_n693, mult_46_n692, mult_46_n691,
         mult_46_n690, mult_46_n689, mult_46_n688, mult_46_n687, mult_46_n686,
         mult_46_n685, mult_46_n684, mult_46_n683, mult_46_n682, mult_46_n681,
         mult_46_n680, mult_46_n679, mult_46_n678, mult_46_n677, mult_46_n676,
         mult_46_n675, mult_46_n674, mult_46_n673, mult_46_n672, mult_46_n671,
         mult_46_n670, mult_46_n669, mult_46_n668, mult_46_n667, mult_46_n666,
         mult_46_n665, mult_46_n664, mult_46_n663, mult_46_n662, mult_46_n661,
         mult_46_n660, mult_46_n659, mult_46_n658, mult_46_n657, mult_46_n656,
         mult_46_n655, mult_46_n654, mult_46_n653, mult_46_n652, mult_46_n651,
         mult_46_n650, mult_46_n649, mult_46_n648, mult_46_n647, mult_46_n646,
         mult_46_n645, mult_46_n644, mult_46_n643, mult_46_n642, mult_46_n641,
         mult_46_n640, mult_46_n639, mult_46_n638, mult_46_n637, mult_46_n636,
         mult_46_n635, mult_46_n419, mult_46_n418, mult_46_n417, mult_46_n416,
         mult_46_n415, mult_46_n414, mult_46_n413, mult_46_n412, mult_46_n411,
         mult_46_n410, mult_46_n409, mult_46_n408, mult_46_n406, mult_46_n405,
         mult_46_n404, mult_46_n403, mult_46_n402, mult_46_n401, mult_46_n400,
         mult_46_n399, mult_46_n398, mult_46_n397, mult_46_n396, mult_46_n395,
         mult_46_n394, mult_46_n393, mult_46_n392, mult_46_n391, mult_46_n390,
         mult_46_n389, mult_46_n388, mult_46_n387, mult_46_n386, mult_46_n385,
         mult_46_n384, mult_46_n382, mult_46_n381, mult_46_n380, mult_46_n379,
         mult_46_n378, mult_46_n377, mult_46_n376, mult_46_n375, mult_46_n374,
         mult_46_n373, mult_46_n372, mult_46_n371, mult_46_n370, mult_46_n369,
         mult_46_n368, mult_46_n367, mult_46_n366, mult_46_n365, mult_46_n364,
         mult_46_n363, mult_46_n362, mult_46_n361, mult_46_n360, mult_46_n359,
         mult_46_n358, mult_46_n357, mult_46_n356, mult_46_n355, mult_46_n354,
         mult_46_n353, mult_46_n352, mult_46_n351, mult_46_n350, mult_46_n349,
         mult_46_n348, mult_46_n346, mult_46_n345, mult_46_n344, mult_46_n343,
         mult_46_n342, mult_46_n341, mult_46_n340, mult_46_n339, mult_46_n338,
         mult_46_n337, mult_46_n336, mult_46_n335, mult_46_n334, mult_46_n333,
         mult_46_n332, mult_46_n331, mult_46_n330, mult_46_n329, mult_46_n328,
         mult_46_n327, mult_46_n326, mult_46_n325, mult_46_n321, mult_46_n320,
         mult_46_n319, mult_46_n318, mult_46_n317, mult_46_n316, mult_46_n315,
         mult_46_n314, mult_46_n313, mult_46_n312, mult_46_n311, mult_46_n310,
         mult_46_n309, mult_46_n308, mult_46_n307, mult_46_n306, mult_46_n305,
         mult_46_n304, mult_46_n303, mult_46_n302, mult_46_n301, mult_46_n300,
         mult_46_n299, mult_46_n298, mult_46_n297, mult_46_n296, mult_46_n295,
         mult_46_n294, mult_46_n293, mult_46_n292, mult_46_n291, mult_46_n290,
         mult_46_n289, mult_46_n288, mult_46_n287, mult_46_n286, mult_46_n285,
         mult_46_n284, mult_46_n283, mult_46_n282, mult_46_n281, mult_46_n280,
         mult_46_n279, mult_46_n278, mult_46_n277, mult_46_n276, mult_46_n275,
         mult_46_n274, mult_46_n273, mult_46_n272, mult_46_n271, mult_46_n270,
         mult_46_n269, mult_46_n268, mult_46_n267, mult_46_n266, mult_46_n265,
         mult_46_n264, mult_46_n263, mult_46_n262, mult_46_n261, mult_46_n260,
         mult_46_n259, mult_46_n258, mult_46_n257, mult_46_n256, mult_46_n255,
         mult_46_n254, mult_46_n253, mult_46_n252, mult_46_n251, mult_46_n250,
         mult_46_n249, mult_46_n248, mult_46_n247, mult_46_n246, mult_46_n245,
         mult_46_n244, mult_46_n243, mult_46_n242, mult_46_n241, mult_46_n240,
         mult_46_n239, mult_46_n238, mult_46_n237, mult_46_n236, mult_46_n235,
         mult_46_n234, mult_46_n233, mult_46_n232, mult_46_n231, mult_46_n230,
         mult_46_n229, mult_46_n228, mult_46_n227, mult_46_n226, mult_46_n225,
         mult_46_n224, mult_46_n223, mult_46_n222, mult_46_n221, mult_46_n220,
         mult_46_n219, mult_46_n218, mult_46_n217, mult_46_n216, mult_46_n215,
         mult_46_n214, mult_46_n213, mult_46_n212, mult_46_n211, mult_46_n210,
         mult_46_n209, mult_46_n208, mult_46_n207, mult_46_n206, mult_46_n205,
         mult_46_n204, mult_46_n203, mult_46_n202, mult_46_n201, mult_46_n200,
         mult_46_n199, mult_46_n198, mult_46_n197, mult_46_n196, mult_46_n195,
         mult_46_n194, mult_46_n193, mult_46_n192, mult_46_n191, mult_46_n190,
         mult_46_n189, mult_46_n188, mult_46_n187, mult_46_n186, mult_46_n185,
         mult_46_n184, mult_46_n183, mult_46_n182, mult_46_n181, mult_46_n180,
         mult_46_n179, mult_46_n178, mult_46_n177, mult_46_n176, mult_46_n175,
         mult_46_n174, mult_46_n173, mult_46_n172, mult_46_n171, mult_46_n170,
         mult_46_n169, mult_46_n168, mult_46_n167, mult_46_n166, mult_46_n165,
         mult_46_n164, mult_46_n163, mult_46_n162, mult_46_n149, mult_46_n148,
         mult_46_n147, mult_46_n146, mult_46_n145, mult_46_n144, mult_46_n143,
         mult_46_n142, mult_46_n141, mult_46_n140, mult_46_n139, mult_46_n138,
         mult_46_n137, mult_46_n136, mult_48_n812, mult_48_n811, mult_48_n810,
         mult_48_n809, mult_48_n808, mult_48_n807, mult_48_n806, mult_48_n805,
         mult_48_n804, mult_48_n803, mult_48_n802, mult_48_n801, mult_48_n800,
         mult_48_n799, mult_48_n798, mult_48_n797, mult_48_n796, mult_48_n795,
         mult_48_n794, mult_48_n793, mult_48_n792, mult_48_n791, mult_48_n790,
         mult_48_n789, mult_48_n788, mult_48_n787, mult_48_n786, mult_48_n785,
         mult_48_n784, mult_48_n783, mult_48_n782, mult_48_n781, mult_48_n780,
         mult_48_n779, mult_48_n778, mult_48_n777, mult_48_n776, mult_48_n775,
         mult_48_n774, mult_48_n773, mult_48_n772, mult_48_n771, mult_48_n770,
         mult_48_n769, mult_48_n768, mult_48_n767, mult_48_n766, mult_48_n765,
         mult_48_n764, mult_48_n763, mult_48_n762, mult_48_n761, mult_48_n760,
         mult_48_n759, mult_48_n758, mult_48_n757, mult_48_n756, mult_48_n755,
         mult_48_n754, mult_48_n753, mult_48_n752, mult_48_n751, mult_48_n750,
         mult_48_n749, mult_48_n748, mult_48_n747, mult_48_n746, mult_48_n745,
         mult_48_n744, mult_48_n743, mult_48_n742, mult_48_n741, mult_48_n740,
         mult_48_n739, mult_48_n738, mult_48_n737, mult_48_n736, mult_48_n735,
         mult_48_n734, mult_48_n733, mult_48_n732, mult_48_n731, mult_48_n730,
         mult_48_n729, mult_48_n728, mult_48_n727, mult_48_n726, mult_48_n725,
         mult_48_n724, mult_48_n723, mult_48_n722, mult_48_n721, mult_48_n720,
         mult_48_n719, mult_48_n718, mult_48_n717, mult_48_n716, mult_48_n715,
         mult_48_n714, mult_48_n713, mult_48_n712, mult_48_n711, mult_48_n710,
         mult_48_n709, mult_48_n708, mult_48_n707, mult_48_n706, mult_48_n705,
         mult_48_n704, mult_48_n703, mult_48_n702, mult_48_n701, mult_48_n700,
         mult_48_n699, mult_48_n698, mult_48_n697, mult_48_n696, mult_48_n695,
         mult_48_n694, mult_48_n693, mult_48_n692, mult_48_n691, mult_48_n690,
         mult_48_n689, mult_48_n688, mult_48_n687, mult_48_n686, mult_48_n685,
         mult_48_n684, mult_48_n683, mult_48_n682, mult_48_n681, mult_48_n680,
         mult_48_n679, mult_48_n678, mult_48_n677, mult_48_n676, mult_48_n675,
         mult_48_n674, mult_48_n673, mult_48_n672, mult_48_n671, mult_48_n670,
         mult_48_n669, mult_48_n668, mult_48_n667, mult_48_n666, mult_48_n665,
         mult_48_n664, mult_48_n663, mult_48_n662, mult_48_n661, mult_48_n660,
         mult_48_n659, mult_48_n658, mult_48_n657, mult_48_n656, mult_48_n655,
         mult_48_n654, mult_48_n653, mult_48_n652, mult_48_n651, mult_48_n650,
         mult_48_n649, mult_48_n648, mult_48_n647, mult_48_n646, mult_48_n645,
         mult_48_n644, mult_48_n643, mult_48_n642, mult_48_n641, mult_48_n640,
         mult_48_n639, mult_48_n638, mult_48_n637, mult_48_n636, mult_48_n635,
         mult_48_n419, mult_48_n418, mult_48_n417, mult_48_n416, mult_48_n415,
         mult_48_n414, mult_48_n413, mult_48_n412, mult_48_n411, mult_48_n410,
         mult_48_n409, mult_48_n408, mult_48_n406, mult_48_n405, mult_48_n404,
         mult_48_n403, mult_48_n402, mult_48_n401, mult_48_n400, mult_48_n399,
         mult_48_n398, mult_48_n397, mult_48_n396, mult_48_n395, mult_48_n394,
         mult_48_n393, mult_48_n392, mult_48_n391, mult_48_n390, mult_48_n389,
         mult_48_n388, mult_48_n387, mult_48_n386, mult_48_n385, mult_48_n384,
         mult_48_n382, mult_48_n381, mult_48_n380, mult_48_n379, mult_48_n378,
         mult_48_n377, mult_48_n376, mult_48_n375, mult_48_n374, mult_48_n373,
         mult_48_n372, mult_48_n371, mult_48_n370, mult_48_n369, mult_48_n368,
         mult_48_n367, mult_48_n366, mult_48_n365, mult_48_n364, mult_48_n363,
         mult_48_n362, mult_48_n361, mult_48_n360, mult_48_n359, mult_48_n358,
         mult_48_n357, mult_48_n356, mult_48_n355, mult_48_n354, mult_48_n353,
         mult_48_n352, mult_48_n351, mult_48_n350, mult_48_n349, mult_48_n348,
         mult_48_n346, mult_48_n345, mult_48_n344, mult_48_n343, mult_48_n342,
         mult_48_n341, mult_48_n340, mult_48_n339, mult_48_n338, mult_48_n337,
         mult_48_n336, mult_48_n335, mult_48_n334, mult_48_n333, mult_48_n332,
         mult_48_n331, mult_48_n330, mult_48_n329, mult_48_n328, mult_48_n327,
         mult_48_n326, mult_48_n325, mult_48_n321, mult_48_n320, mult_48_n319,
         mult_48_n318, mult_48_n317, mult_48_n316, mult_48_n315, mult_48_n314,
         mult_48_n313, mult_48_n312, mult_48_n311, mult_48_n310, mult_48_n309,
         mult_48_n308, mult_48_n307, mult_48_n306, mult_48_n305, mult_48_n304,
         mult_48_n303, mult_48_n302, mult_48_n301, mult_48_n300, mult_48_n299,
         mult_48_n298, mult_48_n297, mult_48_n296, mult_48_n295, mult_48_n294,
         mult_48_n293, mult_48_n292, mult_48_n291, mult_48_n290, mult_48_n289,
         mult_48_n288, mult_48_n287, mult_48_n286, mult_48_n285, mult_48_n284,
         mult_48_n283, mult_48_n282, mult_48_n281, mult_48_n280, mult_48_n279,
         mult_48_n278, mult_48_n277, mult_48_n276, mult_48_n275, mult_48_n274,
         mult_48_n273, mult_48_n272, mult_48_n271, mult_48_n270, mult_48_n269,
         mult_48_n268, mult_48_n267, mult_48_n266, mult_48_n265, mult_48_n264,
         mult_48_n263, mult_48_n262, mult_48_n261, mult_48_n260, mult_48_n259,
         mult_48_n258, mult_48_n257, mult_48_n256, mult_48_n255, mult_48_n254,
         mult_48_n253, mult_48_n252, mult_48_n251, mult_48_n250, mult_48_n249,
         mult_48_n248, mult_48_n247, mult_48_n246, mult_48_n245, mult_48_n244,
         mult_48_n243, mult_48_n242, mult_48_n241, mult_48_n240, mult_48_n239,
         mult_48_n238, mult_48_n237, mult_48_n236, mult_48_n235, mult_48_n234,
         mult_48_n233, mult_48_n232, mult_48_n231, mult_48_n230, mult_48_n229,
         mult_48_n228, mult_48_n227, mult_48_n226, mult_48_n225, mult_48_n224,
         mult_48_n223, mult_48_n222, mult_48_n221, mult_48_n220, mult_48_n219,
         mult_48_n218, mult_48_n217, mult_48_n216, mult_48_n215, mult_48_n214,
         mult_48_n213, mult_48_n212, mult_48_n211, mult_48_n210, mult_48_n209,
         mult_48_n208, mult_48_n207, mult_48_n206, mult_48_n205, mult_48_n204,
         mult_48_n203, mult_48_n202, mult_48_n201, mult_48_n200, mult_48_n199,
         mult_48_n198, mult_48_n197, mult_48_n196, mult_48_n195, mult_48_n194,
         mult_48_n193, mult_48_n192, mult_48_n191, mult_48_n190, mult_48_n189,
         mult_48_n188, mult_48_n187, mult_48_n186, mult_48_n185, mult_48_n184,
         mult_48_n183, mult_48_n182, mult_48_n181, mult_48_n180, mult_48_n179,
         mult_48_n178, mult_48_n177, mult_48_n176, mult_48_n175, mult_48_n174,
         mult_48_n173, mult_48_n172, mult_48_n171, mult_48_n170, mult_48_n169,
         mult_48_n168, mult_48_n167, mult_48_n166, mult_48_n165, mult_48_n164,
         mult_48_n163, mult_48_n162, mult_48_n149, mult_48_n148, mult_48_n147,
         mult_48_n146, mult_48_n145, mult_48_n144, mult_48_n143, mult_48_n142,
         mult_48_n141, mult_48_n140, mult_48_n139, mult_48_n138, mult_48_n137,
         mult_48_n136, sub_1_root_add_0_root_add_58_B_not_0_,
         sub_1_root_add_0_root_add_58_B_not_1_,
         sub_1_root_add_0_root_add_58_B_not_2_,
         sub_1_root_add_0_root_add_58_B_not_3_,
         sub_1_root_add_0_root_add_58_B_not_4_,
         sub_1_root_add_0_root_add_58_B_not_5_,
         sub_1_root_add_0_root_add_58_B_not_6_,
         sub_1_root_add_0_root_add_58_B_not_7_,
         sub_1_root_add_0_root_add_58_B_not_8_,
         sub_1_root_add_0_root_add_58_B_not_9_,
         sub_1_root_add_0_root_add_58_B_not_10_,
         sub_1_root_add_0_root_add_58_B_not_11_,
         sub_1_root_add_0_root_add_58_B_not_12_,
         sub_1_root_add_0_root_add_58_B_not_13_,
         sub_1_root_add_0_root_add_58_carry_1_,
         sub_1_root_add_0_root_add_58_carry_2_,
         sub_1_root_add_0_root_add_58_carry_3_,
         sub_1_root_add_0_root_add_58_carry_4_,
         sub_1_root_add_0_root_add_58_carry_5_,
         sub_1_root_add_0_root_add_58_carry_6_,
         sub_1_root_add_0_root_add_58_carry_7_,
         sub_1_root_add_0_root_add_58_carry_8_,
         sub_1_root_add_0_root_add_58_carry_9_,
         sub_1_root_add_0_root_add_58_carry_10_,
         sub_1_root_add_0_root_add_58_carry_11_,
         sub_1_root_add_0_root_add_58_carry_12_,
         sub_1_root_add_0_root_add_58_carry_13_,
         sub_0_root_add_0_root_add_58_B_not_0_,
         sub_0_root_add_0_root_add_58_B_not_1_,
         sub_0_root_add_0_root_add_58_B_not_2_,
         sub_0_root_add_0_root_add_58_B_not_3_,
         sub_0_root_add_0_root_add_58_B_not_4_,
         sub_0_root_add_0_root_add_58_B_not_5_,
         sub_0_root_add_0_root_add_58_B_not_6_,
         sub_0_root_add_0_root_add_58_B_not_7_,
         sub_0_root_add_0_root_add_58_B_not_8_,
         sub_0_root_add_0_root_add_58_B_not_9_,
         sub_0_root_add_0_root_add_58_B_not_10_,
         sub_0_root_add_0_root_add_58_B_not_11_,
         sub_0_root_add_0_root_add_58_B_not_12_,
         sub_0_root_add_0_root_add_58_B_not_13_,
         sub_0_root_add_0_root_add_58_carry_1_,
         sub_0_root_add_0_root_add_58_carry_2_,
         sub_0_root_add_0_root_add_58_carry_3_,
         sub_0_root_add_0_root_add_58_carry_4_,
         sub_0_root_add_0_root_add_58_carry_5_,
         sub_0_root_add_0_root_add_58_carry_6_,
         sub_0_root_add_0_root_add_58_carry_7_,
         sub_0_root_add_0_root_add_58_carry_8_,
         sub_0_root_add_0_root_add_58_carry_9_,
         sub_0_root_add_0_root_add_58_carry_10_,
         sub_0_root_add_0_root_add_58_carry_11_,
         sub_0_root_add_0_root_add_58_carry_12_,
         sub_0_root_add_0_root_add_58_carry_13_;
  wire   [13:0] reg1;
  wire   [13:0] reg2;
  wire   [13:0] w;

  DFFR_X1 VOUT_reg ( .D(n101), .CK(CLK), .RN(RST_n), .Q(VOUT), .QN(n58) );
  DFFR_X1 reg2_reg_11_ ( .D(n113), .CK(CLK), .RN(RST_n), .Q(n168), .QN(n169)
         );
  DFFR_X1 reg2_reg_9_ ( .D(n111), .CK(CLK), .RN(RST_n), .Q(n166), .QN(n167) );
  DFFR_X1 reg2_reg_4_ ( .D(n106), .CK(CLK), .RN(RST_n), .Q(reg2[4]), .QN(n11)
         );
  DFFR_X1 reg2_reg_2_ ( .D(n104), .CK(CLK), .RN(RST_n), .Q(reg2[2]), .QN(n7)
         );
  DFFR_X1 reg2_reg_1_ ( .D(n103), .CK(CLK), .RN(RST_n), .Q(n158), .QN(n159) );
  DFFR_X1 reg2_reg_13_ ( .D(n115), .CK(CLK), .RN(RST_n), .Q(n170), .QN(n171)
         );
  DFFR_X1 reg2_reg_12_ ( .D(n114), .CK(CLK), .RN(RST_n), .Q(reg2[12]), .QN(n27) );
  DFFR_X1 reg2_reg_10_ ( .D(n112), .CK(CLK), .RN(RST_n), .Q(reg2[10]), .QN(n23) );
  DFFR_X1 reg2_reg_8_ ( .D(n110), .CK(CLK), .RN(RST_n), .Q(reg2[8]), .QN(n19)
         );
  DFFR_X1 reg2_reg_7_ ( .D(n109), .CK(CLK), .RN(RST_n), .Q(n164), .QN(n165) );
  DFFR_X1 reg2_reg_6_ ( .D(n108), .CK(CLK), .RN(RST_n), .Q(reg2[6]), .QN(n15)
         );
  DFFR_X1 reg2_reg_5_ ( .D(n107), .CK(CLK), .RN(RST_n), .Q(n162), .QN(n163) );
  DFFR_X1 reg2_reg_3_ ( .D(n105), .CK(CLK), .RN(RST_n), .Q(n160), .QN(n161) );
  DFFR_X1 reg2_reg_0_ ( .D(n102), .CK(CLK), .RN(RST_n), .Q(reg2[0]), .QN(n3)
         );
  DFFR_X1 xin_reg_1_ ( .D(n131), .CK(CLK), .RN(RST_n), .Q(fb_1_) );
  DFFR_X1 xin_reg_0_ ( .D(n130), .CK(CLK), .RN(RST_n), .Q(fb_0_) );
  DFFR_X1 xin_reg_13_ ( .D(n143), .CK(CLK), .RN(RST_n), .Q(fb_13_) );
  DFFR_X1 xin_reg_12_ ( .D(n142), .CK(CLK), .RN(RST_n), .Q(fb_12_) );
  DFFR_X1 xin_reg_11_ ( .D(n141), .CK(CLK), .RN(RST_n), .Q(fb_11_) );
  DFFR_X1 xin_reg_10_ ( .D(n140), .CK(CLK), .RN(RST_n), .Q(fb_10_) );
  DFFR_X1 xin_reg_9_ ( .D(n139), .CK(CLK), .RN(RST_n), .Q(fb_9_) );
  DFFR_X1 xin_reg_8_ ( .D(n138), .CK(CLK), .RN(RST_n), .Q(fb_8_) );
  DFFR_X1 xin_reg_7_ ( .D(n137), .CK(CLK), .RN(RST_n), .Q(fb_7_) );
  DFFR_X1 xin_reg_6_ ( .D(n136), .CK(CLK), .RN(RST_n), .Q(fb_6_) );
  DFFR_X1 xin_reg_5_ ( .D(n135), .CK(CLK), .RN(RST_n), .Q(fb_5_) );
  DFFR_X1 xin_reg_4_ ( .D(n134), .CK(CLK), .RN(RST_n), .Q(fb_4_) );
  DFFR_X1 xin_reg_3_ ( .D(n133), .CK(CLK), .RN(RST_n), .Q(fb_3_) );
  DFFR_X1 xin_reg_2_ ( .D(n132), .CK(CLK), .RN(RST_n), .Q(fb_2_) );
  DFFR_X1 reg1_reg_0_ ( .D(n116), .CK(CLK), .RN(RST_n), .Q(reg1[0]), .QN(n2)
         );
  DFFR_X1 reg1_reg_2_ ( .D(n118), .CK(CLK), .RN(RST_n), .Q(reg1[2]), .QN(n6)
         );
  DFFR_X1 reg1_reg_1_ ( .D(n117), .CK(CLK), .RN(RST_n), .Q(n172), .QN(n173) );
  DFFR_X1 reg1_reg_4_ ( .D(n120), .CK(CLK), .RN(RST_n), .Q(reg1[4]), .QN(n10)
         );
  DFFR_X1 reg1_reg_3_ ( .D(n119), .CK(CLK), .RN(RST_n), .Q(n174), .QN(n175) );
  DFFR_X1 reg1_reg_6_ ( .D(n122), .CK(CLK), .RN(RST_n), .Q(reg1[6]), .QN(n14)
         );
  DFFR_X1 reg1_reg_5_ ( .D(n121), .CK(CLK), .RN(RST_n), .Q(n176), .QN(n177) );
  DFFR_X1 reg1_reg_8_ ( .D(n124), .CK(CLK), .RN(RST_n), .Q(reg1[8]), .QN(n18)
         );
  DFFR_X1 reg1_reg_7_ ( .D(n123), .CK(CLK), .RN(RST_n), .Q(n178), .QN(n179) );
  DFFR_X1 reg1_reg_10_ ( .D(n126), .CK(CLK), .RN(RST_n), .Q(reg1[10]), .QN(n22) );
  DFFR_X1 reg1_reg_9_ ( .D(n125), .CK(CLK), .RN(RST_n), .Q(n180), .QN(n181) );
  DFFR_X1 reg1_reg_12_ ( .D(n128), .CK(CLK), .RN(RST_n), .Q(reg1[12]), .QN(n26) );
  DFFR_X1 reg1_reg_11_ ( .D(n127), .CK(CLK), .RN(RST_n), .Q(n182), .QN(n183)
         );
  DFFR_X1 reg1_reg_13_ ( .D(n129), .CK(CLK), .RN(RST_n), .Q(n184), .QN(n185)
         );
  INV_X1 U103 ( .A(n204), .ZN(n191) );
  INV_X1 U104 ( .A(n203), .ZN(n189) );
  INV_X1 U105 ( .A(n204), .ZN(n192) );
  INV_X1 U106 ( .A(n203), .ZN(n190) );
  OAI21_X1 U107 ( .B1(n192), .B2(n179), .A(n37), .ZN(n123) );
  NAND2_X1 U108 ( .A1(w[7]), .A2(n191), .ZN(n37) );
  OAI21_X1 U109 ( .B1(n192), .B2(n18), .A(n38), .ZN(n124) );
  NAND2_X1 U110 ( .A1(w[8]), .A2(n191), .ZN(n38) );
  OAI21_X1 U111 ( .B1(n192), .B2(n181), .A(n39), .ZN(n125) );
  NAND2_X1 U112 ( .A1(w[9]), .A2(n190), .ZN(n39) );
  OAI21_X1 U113 ( .B1(n192), .B2(n22), .A(n40), .ZN(n126) );
  NAND2_X1 U114 ( .A1(w[10]), .A2(n190), .ZN(n40) );
  OAI21_X1 U115 ( .B1(n192), .B2(n183), .A(n41), .ZN(n127) );
  NAND2_X1 U116 ( .A1(w[11]), .A2(n190), .ZN(n41) );
  OAI21_X1 U117 ( .B1(n192), .B2(n26), .A(n42), .ZN(n128) );
  NAND2_X1 U118 ( .A1(w[12]), .A2(n190), .ZN(n42) );
  OAI21_X1 U119 ( .B1(n193), .B2(n177), .A(n35), .ZN(n121) );
  NAND2_X1 U120 ( .A1(w[5]), .A2(n191), .ZN(n35) );
  OAI21_X1 U121 ( .B1(n193), .B2(n14), .A(n36), .ZN(n122) );
  NAND2_X1 U122 ( .A1(w[6]), .A2(n191), .ZN(n36) );
  OAI21_X1 U123 ( .B1(n193), .B2(n185), .A(n43), .ZN(n129) );
  NAND2_X1 U124 ( .A1(w[13]), .A2(n190), .ZN(n43) );
  OAI21_X1 U125 ( .B1(n192), .B2(n173), .A(n31), .ZN(n117) );
  NAND2_X1 U126 ( .A1(w[1]), .A2(n190), .ZN(n31) );
  OAI21_X1 U127 ( .B1(n192), .B2(n10), .A(n34), .ZN(n120) );
  NAND2_X1 U128 ( .A1(w[4]), .A2(n190), .ZN(n34) );
  OAI21_X1 U129 ( .B1(n193), .B2(n2), .A(n30), .ZN(n116) );
  NAND2_X1 U130 ( .A1(w[0]), .A2(n190), .ZN(n30) );
  OAI21_X1 U131 ( .B1(n193), .B2(n6), .A(n32), .ZN(n118) );
  NAND2_X1 U132 ( .A1(w[2]), .A2(n190), .ZN(n32) );
  OAI21_X1 U133 ( .B1(n193), .B2(n175), .A(n33), .ZN(n119) );
  NAND2_X1 U134 ( .A1(w[3]), .A2(n190), .ZN(n33) );
  OAI22_X1 U135 ( .A1(n202), .A2(n175), .B1(n191), .B2(n161), .ZN(n105) );
  OAI22_X1 U136 ( .A1(n201), .A2(n177), .B1(n191), .B2(n163), .ZN(n107) );
  OAI22_X1 U137 ( .A1(n200), .A2(n179), .B1(n191), .B2(n165), .ZN(n109) );
  OAI22_X1 U138 ( .A1(n202), .A2(n185), .B1(n191), .B2(n171), .ZN(n115) );
  OAI22_X1 U139 ( .A1(n200), .A2(n173), .B1(n192), .B2(n159), .ZN(n103) );
  OAI22_X1 U140 ( .A1(n199), .A2(n181), .B1(n192), .B2(n167), .ZN(n111) );
  OAI22_X1 U141 ( .A1(n199), .A2(n183), .B1(n192), .B2(n169), .ZN(n113) );
  OAI22_X1 U142 ( .A1(n203), .A2(n2), .B1(n191), .B2(n3), .ZN(n102) );
  OAI22_X1 U143 ( .A1(n201), .A2(n14), .B1(n191), .B2(n15), .ZN(n108) );
  OAI22_X1 U144 ( .A1(n200), .A2(n18), .B1(n191), .B2(n19), .ZN(n110) );
  OAI22_X1 U145 ( .A1(n198), .A2(n22), .B1(n191), .B2(n23), .ZN(n112) );
  OAI22_X1 U146 ( .A1(n198), .A2(n26), .B1(n191), .B2(n27), .ZN(n114) );
  OAI22_X1 U147 ( .A1(n198), .A2(n6), .B1(n192), .B2(n7), .ZN(n104) );
  OAI22_X1 U148 ( .A1(n202), .A2(n10), .B1(n192), .B2(n11), .ZN(n106) );
  BUF_X1 U149 ( .A(VIN), .Z(n186) );
  BUF_X1 U150 ( .A(VIN), .Z(n187) );
  BUF_X1 U151 ( .A(VIN), .Z(n188) );
  NAND2_X1 U152 ( .A1(n58), .A2(n201), .ZN(n101) );
  INV_X1 U153 ( .A(n46), .ZN(n132) );
  AOI22_X1 U154 ( .A1(DIN[2]), .A2(n189), .B1(fb_2_), .B2(n197), .ZN(n46) );
  INV_X1 U155 ( .A(n47), .ZN(n133) );
  AOI22_X1 U156 ( .A1(DIN[3]), .A2(n189), .B1(fb_3_), .B2(n197), .ZN(n47) );
  INV_X1 U157 ( .A(n48), .ZN(n134) );
  AOI22_X1 U158 ( .A1(DIN[4]), .A2(n189), .B1(fb_4_), .B2(n196), .ZN(n48) );
  INV_X1 U159 ( .A(n49), .ZN(n135) );
  AOI22_X1 U160 ( .A1(DIN[5]), .A2(n189), .B1(fb_5_), .B2(n196), .ZN(n49) );
  INV_X1 U161 ( .A(n50), .ZN(n136) );
  AOI22_X1 U162 ( .A1(DIN[6]), .A2(n189), .B1(fb_6_), .B2(n196), .ZN(n50) );
  INV_X1 U163 ( .A(n51), .ZN(n137) );
  AOI22_X1 U164 ( .A1(DIN[7]), .A2(n189), .B1(fb_7_), .B2(n197), .ZN(n51) );
  INV_X1 U165 ( .A(n52), .ZN(n138) );
  AOI22_X1 U166 ( .A1(DIN[8]), .A2(n189), .B1(fb_8_), .B2(n195), .ZN(n52) );
  INV_X1 U167 ( .A(n53), .ZN(n139) );
  AOI22_X1 U168 ( .A1(DIN[9]), .A2(n189), .B1(fb_9_), .B2(n195), .ZN(n53) );
  INV_X1 U169 ( .A(n54), .ZN(n140) );
  AOI22_X1 U170 ( .A1(DIN[10]), .A2(n189), .B1(fb_10_), .B2(n194), .ZN(n54) );
  INV_X1 U171 ( .A(n55), .ZN(n141) );
  AOI22_X1 U172 ( .A1(DIN[11]), .A2(n189), .B1(fb_11_), .B2(n194), .ZN(n55) );
  INV_X1 U173 ( .A(n56), .ZN(n142) );
  AOI22_X1 U174 ( .A1(DIN[12]), .A2(n189), .B1(fb_12_), .B2(n196), .ZN(n56) );
  INV_X1 U175 ( .A(n57), .ZN(n143) );
  AOI22_X1 U176 ( .A1(DIN[13]), .A2(n189), .B1(fb_13_), .B2(n194), .ZN(n57) );
  INV_X1 U177 ( .A(n44), .ZN(n130) );
  AOI22_X1 U178 ( .A1(DIN[0]), .A2(n190), .B1(fb_0_), .B2(n195), .ZN(n44) );
  INV_X1 U179 ( .A(n45), .ZN(n131) );
  AOI22_X1 U180 ( .A1(DIN[1]), .A2(n190), .B1(fb_1_), .B2(n194), .ZN(n45) );
  INV_X1 U181 ( .A(n204), .ZN(n193) );
  INV_X1 U182 ( .A(n186), .ZN(n194) );
  INV_X1 U183 ( .A(n186), .ZN(n195) );
  INV_X1 U184 ( .A(n186), .ZN(n196) );
  INV_X1 U185 ( .A(n186), .ZN(n197) );
  INV_X1 U186 ( .A(n187), .ZN(n198) );
  INV_X1 U187 ( .A(n187), .ZN(n199) );
  INV_X1 U188 ( .A(n187), .ZN(n200) );
  INV_X1 U189 ( .A(n187), .ZN(n201) );
  INV_X1 U190 ( .A(n187), .ZN(n202) );
  INV_X1 U191 ( .A(n188), .ZN(n203) );
  INV_X1 U192 ( .A(n188), .ZN(n204) );
  XOR2_X1 mult_50_U691 ( .A(reg1[2]), .B(n172), .Z(mult_50_n798) );
  NOR2_X1 mult_50_U690 ( .A1(mult_50_n635), .A2(B1[1]), .ZN(mult_50_n803) );
  INV_X1 mult_50_U689 ( .A(mult_50_n803), .ZN(mult_50_n805) );
  NAND2_X1 mult_50_U688 ( .A1(n172), .A2(mult_50_n650), .ZN(mult_50_n648) );
  XNOR2_X1 mult_50_U687 ( .A(B1[2]), .B(n172), .ZN(mult_50_n647) );
  OAI22_X1 mult_50_U686 ( .A1(mult_50_n805), .A2(mult_50_n648), .B1(
        mult_50_n647), .B2(mult_50_n650), .ZN(mult_50_n804) );
  NAND2_X1 mult_50_U685 ( .A1(mult_50_n798), .A2(mult_50_n804), .ZN(
        mult_50_n801) );
  NAND2_X1 mult_50_U684 ( .A1(mult_50_n803), .A2(mult_50_n804), .ZN(
        mult_50_n802) );
  INV_X1 mult_50_U683 ( .A(B1[0]), .ZN(mult_50_n679) );
  MUX2_X1 mult_50_U682 ( .A(mult_50_n801), .B(mult_50_n802), .S(mult_50_n679), 
        .Z(mult_50_n800) );
  INV_X1 mult_50_U681 ( .A(mult_50_n800), .ZN(mult_50_n795) );
  XNOR2_X1 mult_50_U680 ( .A(mult_50_n636), .B(reg1[2]), .ZN(mult_50_n799) );
  NAND2_X1 mult_50_U679 ( .A1(mult_50_n664), .A2(mult_50_n799), .ZN(
        mult_50_n663) );
  NAND3_X1 mult_50_U678 ( .A1(mult_50_n798), .A2(mult_50_n679), .A3(n174), 
        .ZN(mult_50_n797) );
  OAI21_X1 mult_50_U677 ( .B1(mult_50_n636), .B2(mult_50_n663), .A(
        mult_50_n797), .ZN(mult_50_n796) );
  AOI222_X1 mult_50_U676 ( .A1(mult_50_n795), .A2(mult_50_n316), .B1(
        mult_50_n796), .B2(mult_50_n795), .C1(mult_50_n796), .C2(mult_50_n316), 
        .ZN(mult_50_n794) );
  INV_X1 mult_50_U675 ( .A(mult_50_n794), .ZN(mult_50_n793) );
  AOI222_X1 mult_50_U674 ( .A1(mult_50_n793), .A2(mult_50_n314), .B1(
        mult_50_n793), .B2(mult_50_n315), .C1(mult_50_n315), .C2(mult_50_n314), 
        .ZN(mult_50_n792) );
  INV_X1 mult_50_U673 ( .A(mult_50_n792), .ZN(mult_50_n791) );
  AOI222_X1 mult_50_U672 ( .A1(mult_50_n791), .A2(mult_50_n310), .B1(
        mult_50_n791), .B2(mult_50_n313), .C1(mult_50_n313), .C2(mult_50_n310), 
        .ZN(mult_50_n790) );
  INV_X1 mult_50_U671 ( .A(mult_50_n790), .ZN(mult_50_n789) );
  AOI222_X1 mult_50_U670 ( .A1(mult_50_n789), .A2(mult_50_n306), .B1(
        mult_50_n789), .B2(mult_50_n309), .C1(mult_50_n309), .C2(mult_50_n306), 
        .ZN(mult_50_n788) );
  INV_X1 mult_50_U669 ( .A(mult_50_n788), .ZN(mult_50_n787) );
  AOI222_X1 mult_50_U668 ( .A1(mult_50_n787), .A2(mult_50_n300), .B1(
        mult_50_n787), .B2(mult_50_n305), .C1(mult_50_n305), .C2(mult_50_n300), 
        .ZN(mult_50_n786) );
  INV_X1 mult_50_U667 ( .A(mult_50_n786), .ZN(mult_50_n785) );
  AOI222_X1 mult_50_U666 ( .A1(mult_50_n785), .A2(mult_50_n294), .B1(
        mult_50_n785), .B2(mult_50_n299), .C1(mult_50_n299), .C2(mult_50_n294), 
        .ZN(mult_50_n784) );
  INV_X1 mult_50_U665 ( .A(mult_50_n784), .ZN(mult_50_n783) );
  AOI222_X1 mult_50_U664 ( .A1(mult_50_n783), .A2(mult_50_n286), .B1(
        mult_50_n783), .B2(mult_50_n293), .C1(mult_50_n293), .C2(mult_50_n286), 
        .ZN(mult_50_n780) );
  INV_X1 mult_50_U663 ( .A(mult_50_n278), .ZN(mult_50_n781) );
  INV_X1 mult_50_U662 ( .A(mult_50_n285), .ZN(mult_50_n782) );
  OAI222_X1 mult_50_U661 ( .A1(mult_50_n780), .A2(mult_50_n781), .B1(
        mult_50_n780), .B2(mult_50_n782), .C1(mult_50_n782), .C2(mult_50_n781), 
        .ZN(mult_50_n779) );
  AOI222_X1 mult_50_U660 ( .A1(mult_50_n779), .A2(mult_50_n268), .B1(
        mult_50_n779), .B2(mult_50_n277), .C1(mult_50_n277), .C2(mult_50_n268), 
        .ZN(mult_50_n776) );
  INV_X1 mult_50_U659 ( .A(mult_50_n258), .ZN(mult_50_n777) );
  INV_X1 mult_50_U658 ( .A(mult_50_n267), .ZN(mult_50_n778) );
  OAI222_X1 mult_50_U657 ( .A1(mult_50_n776), .A2(mult_50_n777), .B1(
        mult_50_n776), .B2(mult_50_n778), .C1(mult_50_n778), .C2(mult_50_n777), 
        .ZN(mult_50_n149) );
  XOR2_X1 mult_50_U656 ( .A(B1[12]), .B(n184), .Z(mult_50_n763) );
  XNOR2_X1 mult_50_U655 ( .A(mult_50_n641), .B(reg1[12]), .ZN(mult_50_n775) );
  NAND2_X1 mult_50_U654 ( .A1(mult_50_n748), .A2(mult_50_n775), .ZN(
        mult_50_n750) );
  INV_X1 mult_50_U653 ( .A(mult_50_n750), .ZN(mult_50_n644) );
  INV_X1 mult_50_U652 ( .A(mult_50_n748), .ZN(mult_50_n645) );
  XNOR2_X1 mult_50_U651 ( .A(B1[13]), .B(mult_50_n641), .ZN(mult_50_n646) );
  AOI22_X1 mult_50_U650 ( .A1(mult_50_n763), .A2(mult_50_n644), .B1(
        mult_50_n645), .B2(mult_50_n646), .ZN(mult_50_n162) );
  XNOR2_X1 mult_50_U649 ( .A(B1[12]), .B(n182), .ZN(mult_50_n745) );
  XNOR2_X1 mult_50_U648 ( .A(mult_50_n640), .B(reg1[10]), .ZN(mult_50_n774) );
  NAND2_X1 mult_50_U647 ( .A1(mult_50_n731), .A2(mult_50_n774), .ZN(
        mult_50_n733) );
  XNOR2_X1 mult_50_U646 ( .A(B1[13]), .B(n182), .ZN(mult_50_n747) );
  OAI22_X1 mult_50_U645 ( .A1(mult_50_n745), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n747), .ZN(mult_50_n167) );
  INV_X1 mult_50_U644 ( .A(mult_50_n167), .ZN(mult_50_n168) );
  XNOR2_X1 mult_50_U643 ( .A(B1[12]), .B(n180), .ZN(mult_50_n728) );
  XNOR2_X1 mult_50_U642 ( .A(mult_50_n639), .B(reg1[8]), .ZN(mult_50_n773) );
  NAND2_X1 mult_50_U641 ( .A1(mult_50_n714), .A2(mult_50_n773), .ZN(
        mult_50_n716) );
  XNOR2_X1 mult_50_U640 ( .A(B1[13]), .B(n180), .ZN(mult_50_n730) );
  OAI22_X1 mult_50_U639 ( .A1(mult_50_n728), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n730), .ZN(mult_50_n177) );
  INV_X1 mult_50_U638 ( .A(mult_50_n177), .ZN(mult_50_n178) );
  XNOR2_X1 mult_50_U637 ( .A(B1[12]), .B(n178), .ZN(mult_50_n711) );
  XNOR2_X1 mult_50_U636 ( .A(mult_50_n638), .B(reg1[6]), .ZN(mult_50_n772) );
  NAND2_X1 mult_50_U635 ( .A1(mult_50_n697), .A2(mult_50_n772), .ZN(
        mult_50_n699) );
  XNOR2_X1 mult_50_U634 ( .A(B1[13]), .B(n178), .ZN(mult_50_n713) );
  OAI22_X1 mult_50_U633 ( .A1(mult_50_n711), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n713), .ZN(mult_50_n191) );
  INV_X1 mult_50_U632 ( .A(mult_50_n191), .ZN(mult_50_n192) );
  XNOR2_X1 mult_50_U631 ( .A(B1[12]), .B(n176), .ZN(mult_50_n694) );
  XNOR2_X1 mult_50_U630 ( .A(mult_50_n637), .B(reg1[4]), .ZN(mult_50_n771) );
  NAND2_X1 mult_50_U629 ( .A1(mult_50_n680), .A2(mult_50_n771), .ZN(
        mult_50_n682) );
  XNOR2_X1 mult_50_U628 ( .A(B1[13]), .B(n176), .ZN(mult_50_n696) );
  OAI22_X1 mult_50_U627 ( .A1(mult_50_n694), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n696), .ZN(mult_50_n209) );
  INV_X1 mult_50_U626 ( .A(mult_50_n209), .ZN(mult_50_n210) );
  XNOR2_X1 mult_50_U625 ( .A(B1[12]), .B(n174), .ZN(mult_50_n676) );
  XNOR2_X1 mult_50_U624 ( .A(B1[13]), .B(n174), .ZN(mult_50_n678) );
  OAI22_X1 mult_50_U623 ( .A1(mult_50_n676), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n678), .ZN(mult_50_n231) );
  INV_X1 mult_50_U622 ( .A(mult_50_n231), .ZN(mult_50_n232) );
  XNOR2_X1 mult_50_U621 ( .A(B1[3]), .B(n182), .ZN(mult_50_n736) );
  XNOR2_X1 mult_50_U620 ( .A(B1[4]), .B(n182), .ZN(mult_50_n737) );
  OAI22_X1 mult_50_U619 ( .A1(mult_50_n736), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n737), .ZN(mult_50_n769) );
  XNOR2_X1 mult_50_U618 ( .A(B1[9]), .B(n176), .ZN(mult_50_n691) );
  XNOR2_X1 mult_50_U617 ( .A(B1[10]), .B(n176), .ZN(mult_50_n692) );
  OAI22_X1 mult_50_U616 ( .A1(mult_50_n691), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n692), .ZN(mult_50_n770) );
  OR2_X1 mult_50_U615 ( .A1(mult_50_n769), .A2(mult_50_n770), .ZN(mult_50_n243) );
  XNOR2_X1 mult_50_U614 ( .A(mult_50_n769), .B(mult_50_n770), .ZN(mult_50_n244) );
  NAND3_X1 mult_50_U613 ( .A1(mult_50_n645), .A2(mult_50_n679), .A3(n184), 
        .ZN(mult_50_n768) );
  OAI21_X1 mult_50_U612 ( .B1(mult_50_n641), .B2(mult_50_n750), .A(
        mult_50_n768), .ZN(mult_50_n317) );
  OR3_X1 mult_50_U611 ( .A1(mult_50_n731), .A2(B1[0]), .A3(mult_50_n640), .ZN(
        mult_50_n767) );
  OAI21_X1 mult_50_U610 ( .B1(mult_50_n640), .B2(mult_50_n733), .A(
        mult_50_n767), .ZN(mult_50_n318) );
  OR3_X1 mult_50_U609 ( .A1(mult_50_n714), .A2(B1[0]), .A3(mult_50_n639), .ZN(
        mult_50_n766) );
  OAI21_X1 mult_50_U608 ( .B1(mult_50_n639), .B2(mult_50_n716), .A(
        mult_50_n766), .ZN(mult_50_n319) );
  OR3_X1 mult_50_U607 ( .A1(mult_50_n697), .A2(B1[0]), .A3(mult_50_n638), .ZN(
        mult_50_n765) );
  OAI21_X1 mult_50_U606 ( .B1(mult_50_n638), .B2(mult_50_n699), .A(
        mult_50_n765), .ZN(mult_50_n320) );
  OR3_X1 mult_50_U605 ( .A1(mult_50_n680), .A2(B1[0]), .A3(mult_50_n637), .ZN(
        mult_50_n764) );
  OAI21_X1 mult_50_U604 ( .B1(mult_50_n637), .B2(mult_50_n682), .A(
        mult_50_n764), .ZN(mult_50_n321) );
  XNOR2_X1 mult_50_U603 ( .A(B1[11]), .B(n184), .ZN(mult_50_n761) );
  INV_X1 mult_50_U602 ( .A(mult_50_n763), .ZN(mult_50_n762) );
  OAI22_X1 mult_50_U601 ( .A1(mult_50_n761), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n762), .ZN(mult_50_n325) );
  XNOR2_X1 mult_50_U600 ( .A(B1[10]), .B(n184), .ZN(mult_50_n760) );
  OAI22_X1 mult_50_U599 ( .A1(mult_50_n760), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n761), .ZN(mult_50_n326) );
  XNOR2_X1 mult_50_U598 ( .A(B1[9]), .B(n184), .ZN(mult_50_n759) );
  OAI22_X1 mult_50_U597 ( .A1(mult_50_n759), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n760), .ZN(mult_50_n327) );
  XNOR2_X1 mult_50_U596 ( .A(B1[8]), .B(n184), .ZN(mult_50_n758) );
  OAI22_X1 mult_50_U595 ( .A1(mult_50_n758), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n759), .ZN(mult_50_n328) );
  XNOR2_X1 mult_50_U594 ( .A(B1[7]), .B(n184), .ZN(mult_50_n757) );
  OAI22_X1 mult_50_U593 ( .A1(mult_50_n757), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n758), .ZN(mult_50_n329) );
  XNOR2_X1 mult_50_U592 ( .A(B1[6]), .B(n184), .ZN(mult_50_n756) );
  OAI22_X1 mult_50_U591 ( .A1(mult_50_n756), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n757), .ZN(mult_50_n330) );
  XNOR2_X1 mult_50_U590 ( .A(B1[5]), .B(n184), .ZN(mult_50_n755) );
  OAI22_X1 mult_50_U589 ( .A1(mult_50_n755), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n756), .ZN(mult_50_n331) );
  XNOR2_X1 mult_50_U588 ( .A(B1[4]), .B(n184), .ZN(mult_50_n754) );
  OAI22_X1 mult_50_U587 ( .A1(mult_50_n754), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n755), .ZN(mult_50_n332) );
  XNOR2_X1 mult_50_U586 ( .A(B1[3]), .B(n184), .ZN(mult_50_n753) );
  OAI22_X1 mult_50_U585 ( .A1(mult_50_n753), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n754), .ZN(mult_50_n333) );
  XNOR2_X1 mult_50_U584 ( .A(B1[2]), .B(n184), .ZN(mult_50_n752) );
  OAI22_X1 mult_50_U583 ( .A1(mult_50_n752), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n753), .ZN(mult_50_n334) );
  XNOR2_X1 mult_50_U582 ( .A(B1[1]), .B(n184), .ZN(mult_50_n751) );
  OAI22_X1 mult_50_U581 ( .A1(mult_50_n751), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n752), .ZN(mult_50_n335) );
  XNOR2_X1 mult_50_U580 ( .A(n184), .B(B1[0]), .ZN(mult_50_n749) );
  OAI22_X1 mult_50_U579 ( .A1(mult_50_n749), .A2(mult_50_n750), .B1(
        mult_50_n748), .B2(mult_50_n751), .ZN(mult_50_n336) );
  NOR2_X1 mult_50_U578 ( .A1(mult_50_n679), .A2(mult_50_n748), .ZN(
        mult_50_n337) );
  AOI21_X1 mult_50_U577 ( .B1(mult_50_n733), .B2(mult_50_n731), .A(
        mult_50_n747), .ZN(mult_50_n746) );
  INV_X1 mult_50_U576 ( .A(mult_50_n746), .ZN(mult_50_n338) );
  XNOR2_X1 mult_50_U575 ( .A(B1[11]), .B(n182), .ZN(mult_50_n744) );
  OAI22_X1 mult_50_U574 ( .A1(mult_50_n744), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n745), .ZN(mult_50_n339) );
  XNOR2_X1 mult_50_U573 ( .A(B1[10]), .B(n182), .ZN(mult_50_n743) );
  OAI22_X1 mult_50_U572 ( .A1(mult_50_n743), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n744), .ZN(mult_50_n340) );
  XNOR2_X1 mult_50_U571 ( .A(B1[9]), .B(n182), .ZN(mult_50_n742) );
  OAI22_X1 mult_50_U570 ( .A1(mult_50_n742), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n743), .ZN(mult_50_n341) );
  XNOR2_X1 mult_50_U569 ( .A(B1[8]), .B(n182), .ZN(mult_50_n741) );
  OAI22_X1 mult_50_U568 ( .A1(mult_50_n741), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n742), .ZN(mult_50_n342) );
  XNOR2_X1 mult_50_U567 ( .A(B1[7]), .B(n182), .ZN(mult_50_n740) );
  OAI22_X1 mult_50_U566 ( .A1(mult_50_n740), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n741), .ZN(mult_50_n343) );
  XNOR2_X1 mult_50_U565 ( .A(B1[6]), .B(n182), .ZN(mult_50_n739) );
  OAI22_X1 mult_50_U564 ( .A1(mult_50_n739), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n740), .ZN(mult_50_n344) );
  XNOR2_X1 mult_50_U563 ( .A(B1[5]), .B(n182), .ZN(mult_50_n738) );
  OAI22_X1 mult_50_U562 ( .A1(mult_50_n738), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n739), .ZN(mult_50_n345) );
  OAI22_X1 mult_50_U561 ( .A1(mult_50_n737), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n738), .ZN(mult_50_n346) );
  XNOR2_X1 mult_50_U560 ( .A(B1[2]), .B(n182), .ZN(mult_50_n735) );
  OAI22_X1 mult_50_U559 ( .A1(mult_50_n735), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n736), .ZN(mult_50_n348) );
  XNOR2_X1 mult_50_U558 ( .A(B1[1]), .B(n182), .ZN(mult_50_n734) );
  OAI22_X1 mult_50_U557 ( .A1(mult_50_n734), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n735), .ZN(mult_50_n349) );
  XNOR2_X1 mult_50_U556 ( .A(n182), .B(B1[0]), .ZN(mult_50_n732) );
  OAI22_X1 mult_50_U555 ( .A1(mult_50_n732), .A2(mult_50_n733), .B1(
        mult_50_n731), .B2(mult_50_n734), .ZN(mult_50_n350) );
  NOR2_X1 mult_50_U554 ( .A1(mult_50_n679), .A2(mult_50_n731), .ZN(
        mult_50_n351) );
  AOI21_X1 mult_50_U553 ( .B1(mult_50_n716), .B2(mult_50_n714), .A(
        mult_50_n730), .ZN(mult_50_n729) );
  INV_X1 mult_50_U552 ( .A(mult_50_n729), .ZN(mult_50_n352) );
  XNOR2_X1 mult_50_U551 ( .A(B1[11]), .B(n180), .ZN(mult_50_n727) );
  OAI22_X1 mult_50_U550 ( .A1(mult_50_n727), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n728), .ZN(mult_50_n353) );
  XNOR2_X1 mult_50_U549 ( .A(B1[10]), .B(n180), .ZN(mult_50_n726) );
  OAI22_X1 mult_50_U548 ( .A1(mult_50_n726), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n727), .ZN(mult_50_n354) );
  XNOR2_X1 mult_50_U547 ( .A(B1[9]), .B(n180), .ZN(mult_50_n725) );
  OAI22_X1 mult_50_U546 ( .A1(mult_50_n725), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n726), .ZN(mult_50_n355) );
  XNOR2_X1 mult_50_U545 ( .A(B1[8]), .B(n180), .ZN(mult_50_n724) );
  OAI22_X1 mult_50_U544 ( .A1(mult_50_n724), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n725), .ZN(mult_50_n356) );
  XNOR2_X1 mult_50_U543 ( .A(B1[7]), .B(n180), .ZN(mult_50_n723) );
  OAI22_X1 mult_50_U542 ( .A1(mult_50_n723), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n724), .ZN(mult_50_n357) );
  XNOR2_X1 mult_50_U541 ( .A(B1[6]), .B(n180), .ZN(mult_50_n722) );
  OAI22_X1 mult_50_U540 ( .A1(mult_50_n722), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n723), .ZN(mult_50_n358) );
  XNOR2_X1 mult_50_U539 ( .A(B1[5]), .B(n180), .ZN(mult_50_n721) );
  OAI22_X1 mult_50_U538 ( .A1(mult_50_n721), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n722), .ZN(mult_50_n359) );
  XNOR2_X1 mult_50_U537 ( .A(B1[4]), .B(n180), .ZN(mult_50_n720) );
  OAI22_X1 mult_50_U536 ( .A1(mult_50_n720), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n721), .ZN(mult_50_n360) );
  XNOR2_X1 mult_50_U535 ( .A(B1[3]), .B(n180), .ZN(mult_50_n719) );
  OAI22_X1 mult_50_U534 ( .A1(mult_50_n719), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n720), .ZN(mult_50_n361) );
  XNOR2_X1 mult_50_U533 ( .A(B1[2]), .B(n180), .ZN(mult_50_n718) );
  OAI22_X1 mult_50_U532 ( .A1(mult_50_n718), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n719), .ZN(mult_50_n362) );
  XNOR2_X1 mult_50_U531 ( .A(B1[1]), .B(n180), .ZN(mult_50_n717) );
  OAI22_X1 mult_50_U530 ( .A1(mult_50_n717), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n718), .ZN(mult_50_n363) );
  XNOR2_X1 mult_50_U529 ( .A(n180), .B(B1[0]), .ZN(mult_50_n715) );
  OAI22_X1 mult_50_U528 ( .A1(mult_50_n715), .A2(mult_50_n716), .B1(
        mult_50_n714), .B2(mult_50_n717), .ZN(mult_50_n364) );
  NOR2_X1 mult_50_U527 ( .A1(mult_50_n679), .A2(mult_50_n714), .ZN(
        mult_50_n365) );
  AOI21_X1 mult_50_U526 ( .B1(mult_50_n699), .B2(mult_50_n697), .A(
        mult_50_n713), .ZN(mult_50_n712) );
  INV_X1 mult_50_U525 ( .A(mult_50_n712), .ZN(mult_50_n366) );
  XNOR2_X1 mult_50_U524 ( .A(B1[11]), .B(n178), .ZN(mult_50_n710) );
  OAI22_X1 mult_50_U523 ( .A1(mult_50_n710), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n711), .ZN(mult_50_n367) );
  XNOR2_X1 mult_50_U522 ( .A(B1[10]), .B(n178), .ZN(mult_50_n709) );
  OAI22_X1 mult_50_U521 ( .A1(mult_50_n709), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n710), .ZN(mult_50_n368) );
  XNOR2_X1 mult_50_U520 ( .A(B1[9]), .B(n178), .ZN(mult_50_n708) );
  OAI22_X1 mult_50_U519 ( .A1(mult_50_n708), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n709), .ZN(mult_50_n369) );
  XNOR2_X1 mult_50_U518 ( .A(B1[8]), .B(n178), .ZN(mult_50_n707) );
  OAI22_X1 mult_50_U517 ( .A1(mult_50_n707), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n708), .ZN(mult_50_n370) );
  XNOR2_X1 mult_50_U516 ( .A(B1[7]), .B(n178), .ZN(mult_50_n706) );
  OAI22_X1 mult_50_U515 ( .A1(mult_50_n706), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n707), .ZN(mult_50_n371) );
  XNOR2_X1 mult_50_U514 ( .A(B1[6]), .B(n178), .ZN(mult_50_n705) );
  OAI22_X1 mult_50_U513 ( .A1(mult_50_n705), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n706), .ZN(mult_50_n372) );
  XNOR2_X1 mult_50_U512 ( .A(B1[5]), .B(n178), .ZN(mult_50_n704) );
  OAI22_X1 mult_50_U511 ( .A1(mult_50_n704), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n705), .ZN(mult_50_n373) );
  XNOR2_X1 mult_50_U510 ( .A(B1[4]), .B(n178), .ZN(mult_50_n703) );
  OAI22_X1 mult_50_U509 ( .A1(mult_50_n703), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n704), .ZN(mult_50_n374) );
  XNOR2_X1 mult_50_U508 ( .A(B1[3]), .B(n178), .ZN(mult_50_n702) );
  OAI22_X1 mult_50_U507 ( .A1(mult_50_n702), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n703), .ZN(mult_50_n375) );
  XNOR2_X1 mult_50_U506 ( .A(B1[2]), .B(n178), .ZN(mult_50_n701) );
  OAI22_X1 mult_50_U505 ( .A1(mult_50_n701), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n702), .ZN(mult_50_n376) );
  XNOR2_X1 mult_50_U504 ( .A(B1[1]), .B(n178), .ZN(mult_50_n700) );
  OAI22_X1 mult_50_U503 ( .A1(mult_50_n700), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n701), .ZN(mult_50_n377) );
  XNOR2_X1 mult_50_U502 ( .A(n178), .B(B1[0]), .ZN(mult_50_n698) );
  OAI22_X1 mult_50_U501 ( .A1(mult_50_n698), .A2(mult_50_n699), .B1(
        mult_50_n697), .B2(mult_50_n700), .ZN(mult_50_n378) );
  NOR2_X1 mult_50_U500 ( .A1(mult_50_n679), .A2(mult_50_n697), .ZN(
        mult_50_n379) );
  AOI21_X1 mult_50_U499 ( .B1(mult_50_n682), .B2(mult_50_n680), .A(
        mult_50_n696), .ZN(mult_50_n695) );
  INV_X1 mult_50_U498 ( .A(mult_50_n695), .ZN(mult_50_n380) );
  XNOR2_X1 mult_50_U497 ( .A(B1[11]), .B(n176), .ZN(mult_50_n693) );
  OAI22_X1 mult_50_U496 ( .A1(mult_50_n693), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n694), .ZN(mult_50_n381) );
  OAI22_X1 mult_50_U495 ( .A1(mult_50_n692), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n693), .ZN(mult_50_n382) );
  XNOR2_X1 mult_50_U494 ( .A(B1[8]), .B(n176), .ZN(mult_50_n690) );
  OAI22_X1 mult_50_U493 ( .A1(mult_50_n690), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n691), .ZN(mult_50_n384) );
  XNOR2_X1 mult_50_U492 ( .A(B1[7]), .B(n176), .ZN(mult_50_n689) );
  OAI22_X1 mult_50_U491 ( .A1(mult_50_n689), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n690), .ZN(mult_50_n385) );
  XNOR2_X1 mult_50_U490 ( .A(B1[6]), .B(n176), .ZN(mult_50_n688) );
  OAI22_X1 mult_50_U489 ( .A1(mult_50_n688), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n689), .ZN(mult_50_n386) );
  XNOR2_X1 mult_50_U488 ( .A(B1[5]), .B(n176), .ZN(mult_50_n687) );
  OAI22_X1 mult_50_U487 ( .A1(mult_50_n687), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n688), .ZN(mult_50_n387) );
  XNOR2_X1 mult_50_U486 ( .A(B1[4]), .B(n176), .ZN(mult_50_n686) );
  OAI22_X1 mult_50_U485 ( .A1(mult_50_n686), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n687), .ZN(mult_50_n388) );
  XNOR2_X1 mult_50_U484 ( .A(B1[3]), .B(n176), .ZN(mult_50_n685) );
  OAI22_X1 mult_50_U483 ( .A1(mult_50_n685), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n686), .ZN(mult_50_n389) );
  XNOR2_X1 mult_50_U482 ( .A(B1[2]), .B(n176), .ZN(mult_50_n684) );
  OAI22_X1 mult_50_U481 ( .A1(mult_50_n684), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n685), .ZN(mult_50_n390) );
  XNOR2_X1 mult_50_U480 ( .A(B1[1]), .B(n176), .ZN(mult_50_n683) );
  OAI22_X1 mult_50_U479 ( .A1(mult_50_n683), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n684), .ZN(mult_50_n391) );
  XNOR2_X1 mult_50_U478 ( .A(n176), .B(B1[0]), .ZN(mult_50_n681) );
  OAI22_X1 mult_50_U477 ( .A1(mult_50_n681), .A2(mult_50_n682), .B1(
        mult_50_n680), .B2(mult_50_n683), .ZN(mult_50_n392) );
  NOR2_X1 mult_50_U476 ( .A1(mult_50_n679), .A2(mult_50_n680), .ZN(
        mult_50_n393) );
  AOI21_X1 mult_50_U475 ( .B1(mult_50_n663), .B2(mult_50_n664), .A(
        mult_50_n678), .ZN(mult_50_n677) );
  INV_X1 mult_50_U474 ( .A(mult_50_n677), .ZN(mult_50_n394) );
  XNOR2_X1 mult_50_U473 ( .A(B1[11]), .B(n174), .ZN(mult_50_n675) );
  OAI22_X1 mult_50_U472 ( .A1(mult_50_n675), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n676), .ZN(mult_50_n395) );
  XNOR2_X1 mult_50_U471 ( .A(B1[10]), .B(n174), .ZN(mult_50_n674) );
  OAI22_X1 mult_50_U470 ( .A1(mult_50_n674), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n675), .ZN(mult_50_n396) );
  XNOR2_X1 mult_50_U469 ( .A(B1[9]), .B(n174), .ZN(mult_50_n673) );
  OAI22_X1 mult_50_U468 ( .A1(mult_50_n673), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n674), .ZN(mult_50_n397) );
  XNOR2_X1 mult_50_U467 ( .A(B1[8]), .B(n174), .ZN(mult_50_n672) );
  OAI22_X1 mult_50_U466 ( .A1(mult_50_n672), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n673), .ZN(mult_50_n398) );
  XNOR2_X1 mult_50_U465 ( .A(B1[7]), .B(n174), .ZN(mult_50_n671) );
  OAI22_X1 mult_50_U464 ( .A1(mult_50_n671), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n672), .ZN(mult_50_n399) );
  XNOR2_X1 mult_50_U463 ( .A(B1[6]), .B(n174), .ZN(mult_50_n670) );
  OAI22_X1 mult_50_U462 ( .A1(mult_50_n670), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n671), .ZN(mult_50_n400) );
  XNOR2_X1 mult_50_U461 ( .A(B1[5]), .B(n174), .ZN(mult_50_n669) );
  OAI22_X1 mult_50_U460 ( .A1(mult_50_n669), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n670), .ZN(mult_50_n401) );
  XNOR2_X1 mult_50_U459 ( .A(B1[4]), .B(n174), .ZN(mult_50_n668) );
  OAI22_X1 mult_50_U458 ( .A1(mult_50_n668), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n669), .ZN(mult_50_n402) );
  XNOR2_X1 mult_50_U457 ( .A(B1[3]), .B(n174), .ZN(mult_50_n667) );
  OAI22_X1 mult_50_U456 ( .A1(mult_50_n667), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n668), .ZN(mult_50_n403) );
  XNOR2_X1 mult_50_U455 ( .A(B1[2]), .B(n174), .ZN(mult_50_n666) );
  OAI22_X1 mult_50_U454 ( .A1(mult_50_n666), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n667), .ZN(mult_50_n404) );
  XNOR2_X1 mult_50_U453 ( .A(B1[1]), .B(n174), .ZN(mult_50_n665) );
  OAI22_X1 mult_50_U452 ( .A1(mult_50_n665), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n666), .ZN(mult_50_n405) );
  XNOR2_X1 mult_50_U451 ( .A(n174), .B(B1[0]), .ZN(mult_50_n662) );
  OAI22_X1 mult_50_U450 ( .A1(mult_50_n662), .A2(mult_50_n663), .B1(
        mult_50_n664), .B2(mult_50_n665), .ZN(mult_50_n406) );
  XOR2_X1 mult_50_U449 ( .A(B1[13]), .B(mult_50_n635), .Z(mult_50_n660) );
  AOI21_X1 mult_50_U448 ( .B1(mult_50_n648), .B2(mult_50_n650), .A(
        mult_50_n660), .ZN(mult_50_n661) );
  INV_X1 mult_50_U447 ( .A(mult_50_n661), .ZN(mult_50_n408) );
  XNOR2_X1 mult_50_U446 ( .A(B1[12]), .B(n172), .ZN(mult_50_n659) );
  OAI22_X1 mult_50_U445 ( .A1(mult_50_n659), .A2(mult_50_n648), .B1(
        mult_50_n660), .B2(mult_50_n650), .ZN(mult_50_n409) );
  XNOR2_X1 mult_50_U444 ( .A(B1[11]), .B(n172), .ZN(mult_50_n658) );
  OAI22_X1 mult_50_U443 ( .A1(mult_50_n658), .A2(mult_50_n648), .B1(
        mult_50_n659), .B2(mult_50_n650), .ZN(mult_50_n410) );
  XNOR2_X1 mult_50_U442 ( .A(B1[10]), .B(n172), .ZN(mult_50_n657) );
  OAI22_X1 mult_50_U441 ( .A1(mult_50_n657), .A2(mult_50_n648), .B1(
        mult_50_n658), .B2(mult_50_n650), .ZN(mult_50_n411) );
  XNOR2_X1 mult_50_U440 ( .A(B1[9]), .B(n172), .ZN(mult_50_n656) );
  OAI22_X1 mult_50_U439 ( .A1(mult_50_n656), .A2(mult_50_n648), .B1(
        mult_50_n657), .B2(mult_50_n650), .ZN(mult_50_n412) );
  XNOR2_X1 mult_50_U438 ( .A(B1[8]), .B(n172), .ZN(mult_50_n655) );
  OAI22_X1 mult_50_U437 ( .A1(mult_50_n655), .A2(mult_50_n648), .B1(
        mult_50_n656), .B2(mult_50_n650), .ZN(mult_50_n413) );
  XNOR2_X1 mult_50_U436 ( .A(B1[7]), .B(n172), .ZN(mult_50_n654) );
  OAI22_X1 mult_50_U435 ( .A1(mult_50_n654), .A2(mult_50_n648), .B1(
        mult_50_n655), .B2(mult_50_n650), .ZN(mult_50_n414) );
  XNOR2_X1 mult_50_U434 ( .A(B1[6]), .B(n172), .ZN(mult_50_n653) );
  OAI22_X1 mult_50_U433 ( .A1(mult_50_n653), .A2(mult_50_n648), .B1(
        mult_50_n654), .B2(mult_50_n650), .ZN(mult_50_n415) );
  XNOR2_X1 mult_50_U432 ( .A(B1[5]), .B(n172), .ZN(mult_50_n652) );
  OAI22_X1 mult_50_U431 ( .A1(mult_50_n652), .A2(mult_50_n648), .B1(
        mult_50_n653), .B2(mult_50_n650), .ZN(mult_50_n416) );
  XNOR2_X1 mult_50_U430 ( .A(B1[4]), .B(n172), .ZN(mult_50_n651) );
  OAI22_X1 mult_50_U429 ( .A1(mult_50_n651), .A2(mult_50_n648), .B1(
        mult_50_n652), .B2(mult_50_n650), .ZN(mult_50_n417) );
  XNOR2_X1 mult_50_U428 ( .A(B1[3]), .B(n172), .ZN(mult_50_n649) );
  OAI22_X1 mult_50_U427 ( .A1(mult_50_n649), .A2(mult_50_n648), .B1(
        mult_50_n651), .B2(mult_50_n650), .ZN(mult_50_n418) );
  OAI22_X1 mult_50_U426 ( .A1(mult_50_n647), .A2(mult_50_n648), .B1(
        mult_50_n649), .B2(mult_50_n650), .ZN(mult_50_n419) );
  OAI21_X1 mult_50_U425 ( .B1(mult_50_n644), .B2(mult_50_n645), .A(
        mult_50_n646), .ZN(mult_50_n643) );
  XOR2_X1 mult_50_U424 ( .A(mult_50_n643), .B(mult_50_n136), .Z(mult_50_n642)
         );
  XNOR2_X1 mult_50_U423 ( .A(mult_50_n162), .B(mult_50_n642), .ZN(temp3_26_)
         );
  INV_X1 mult_50_U422 ( .A(n182), .ZN(mult_50_n640) );
  INV_X1 mult_50_U421 ( .A(n180), .ZN(mult_50_n639) );
  INV_X1 mult_50_U420 ( .A(n178), .ZN(mult_50_n638) );
  INV_X1 mult_50_U419 ( .A(n176), .ZN(mult_50_n637) );
  XOR2_X2 mult_50_U418 ( .A(reg1[12]), .B(mult_50_n640), .Z(mult_50_n748) );
  XOR2_X2 mult_50_U417 ( .A(reg1[10]), .B(mult_50_n639), .Z(mult_50_n731) );
  XOR2_X2 mult_50_U416 ( .A(reg1[8]), .B(mult_50_n638), .Z(mult_50_n714) );
  XOR2_X2 mult_50_U415 ( .A(reg1[6]), .B(mult_50_n637), .Z(mult_50_n697) );
  XOR2_X2 mult_50_U414 ( .A(reg1[4]), .B(mult_50_n636), .Z(mult_50_n680) );
  INV_X1 mult_50_U413 ( .A(reg1[0]), .ZN(mult_50_n650) );
  INV_X1 mult_50_U412 ( .A(mult_50_n798), .ZN(mult_50_n664) );
  INV_X1 mult_50_U411 ( .A(n184), .ZN(mult_50_n641) );
  INV_X1 mult_50_U410 ( .A(n174), .ZN(mult_50_n636) );
  INV_X1 mult_50_U409 ( .A(n172), .ZN(mult_50_n635) );
  HA_X1 mult_50_U145 ( .A(mult_50_n406), .B(mult_50_n419), .CO(mult_50_n315), 
        .S(mult_50_n316) );
  FA_X1 mult_50_U144 ( .A(mult_50_n418), .B(mult_50_n393), .CI(mult_50_n405), 
        .CO(mult_50_n313), .S(mult_50_n314) );
  HA_X1 mult_50_U143 ( .A(mult_50_n321), .B(mult_50_n392), .CO(mult_50_n311), 
        .S(mult_50_n312) );
  FA_X1 mult_50_U142 ( .A(mult_50_n404), .B(mult_50_n417), .CI(mult_50_n312), 
        .CO(mult_50_n309), .S(mult_50_n310) );
  FA_X1 mult_50_U141 ( .A(mult_50_n416), .B(mult_50_n379), .CI(mult_50_n403), 
        .CO(mult_50_n307), .S(mult_50_n308) );
  FA_X1 mult_50_U140 ( .A(mult_50_n311), .B(mult_50_n391), .CI(mult_50_n308), 
        .CO(mult_50_n305), .S(mult_50_n306) );
  HA_X1 mult_50_U139 ( .A(mult_50_n320), .B(mult_50_n378), .CO(mult_50_n303), 
        .S(mult_50_n304) );
  FA_X1 mult_50_U138 ( .A(mult_50_n390), .B(mult_50_n415), .CI(mult_50_n402), 
        .CO(mult_50_n301), .S(mult_50_n302) );
  FA_X1 mult_50_U137 ( .A(mult_50_n307), .B(mult_50_n304), .CI(mult_50_n302), 
        .CO(mult_50_n299), .S(mult_50_n300) );
  FA_X1 mult_50_U136 ( .A(mult_50_n389), .B(mult_50_n365), .CI(mult_50_n414), 
        .CO(mult_50_n297), .S(mult_50_n298) );
  FA_X1 mult_50_U135 ( .A(mult_50_n377), .B(mult_50_n401), .CI(mult_50_n303), 
        .CO(mult_50_n295), .S(mult_50_n296) );
  FA_X1 mult_50_U134 ( .A(mult_50_n298), .B(mult_50_n301), .CI(mult_50_n296), 
        .CO(mult_50_n293), .S(mult_50_n294) );
  HA_X1 mult_50_U133 ( .A(mult_50_n319), .B(mult_50_n364), .CO(mult_50_n291), 
        .S(mult_50_n292) );
  FA_X1 mult_50_U132 ( .A(mult_50_n376), .B(mult_50_n388), .CI(mult_50_n400), 
        .CO(mult_50_n289), .S(mult_50_n290) );
  FA_X1 mult_50_U131 ( .A(mult_50_n292), .B(mult_50_n413), .CI(mult_50_n297), 
        .CO(mult_50_n287), .S(mult_50_n288) );
  FA_X1 mult_50_U130 ( .A(mult_50_n290), .B(mult_50_n295), .CI(mult_50_n288), 
        .CO(mult_50_n285), .S(mult_50_n286) );
  FA_X1 mult_50_U129 ( .A(mult_50_n375), .B(mult_50_n351), .CI(mult_50_n412), 
        .CO(mult_50_n283), .S(mult_50_n284) );
  FA_X1 mult_50_U128 ( .A(mult_50_n363), .B(mult_50_n399), .CI(mult_50_n387), 
        .CO(mult_50_n281), .S(mult_50_n282) );
  FA_X1 mult_50_U127 ( .A(mult_50_n289), .B(mult_50_n291), .CI(mult_50_n284), 
        .CO(mult_50_n279), .S(mult_50_n280) );
  FA_X1 mult_50_U126 ( .A(mult_50_n287), .B(mult_50_n282), .CI(mult_50_n280), 
        .CO(mult_50_n277), .S(mult_50_n278) );
  HA_X1 mult_50_U125 ( .A(mult_50_n318), .B(mult_50_n350), .CO(mult_50_n275), 
        .S(mult_50_n276) );
  FA_X1 mult_50_U124 ( .A(mult_50_n362), .B(mult_50_n386), .CI(mult_50_n411), 
        .CO(mult_50_n273), .S(mult_50_n274) );
  FA_X1 mult_50_U123 ( .A(mult_50_n374), .B(mult_50_n398), .CI(mult_50_n276), 
        .CO(mult_50_n271), .S(mult_50_n272) );
  FA_X1 mult_50_U122 ( .A(mult_50_n281), .B(mult_50_n283), .CI(mult_50_n274), 
        .CO(mult_50_n269), .S(mult_50_n270) );
  FA_X1 mult_50_U121 ( .A(mult_50_n279), .B(mult_50_n272), .CI(mult_50_n270), 
        .CO(mult_50_n267), .S(mult_50_n268) );
  FA_X1 mult_50_U120 ( .A(mult_50_n361), .B(mult_50_n337), .CI(mult_50_n410), 
        .CO(mult_50_n265), .S(mult_50_n266) );
  FA_X1 mult_50_U109 ( .A(mult_50_n349), .B(mult_50_n397), .CI(mult_50_n373), 
        .CO(mult_50_n263), .S(mult_50_n264) );
  FA_X1 mult_50_U108 ( .A(mult_50_n275), .B(mult_50_n385), .CI(mult_50_n273), 
        .CO(mult_50_n261), .S(mult_50_n262) );
  FA_X1 mult_50_U107 ( .A(mult_50_n264), .B(mult_50_n266), .CI(mult_50_n271), 
        .CO(mult_50_n259), .S(mult_50_n260) );
  FA_X1 mult_50_U106 ( .A(mult_50_n262), .B(mult_50_n269), .CI(mult_50_n260), 
        .CO(mult_50_n257), .S(mult_50_n258) );
  HA_X1 mult_50_U105 ( .A(mult_50_n317), .B(mult_50_n336), .CO(mult_50_n255), 
        .S(mult_50_n256) );
  FA_X1 mult_50_U104 ( .A(mult_50_n409), .B(mult_50_n372), .CI(mult_50_n396), 
        .CO(mult_50_n253), .S(mult_50_n254) );
  FA_X1 mult_50_U103 ( .A(mult_50_n348), .B(mult_50_n384), .CI(mult_50_n360), 
        .CO(mult_50_n251), .S(mult_50_n252) );
  FA_X1 mult_50_U102 ( .A(mult_50_n265), .B(mult_50_n256), .CI(mult_50_n263), 
        .CO(mult_50_n249), .S(mult_50_n250) );
  FA_X1 mult_50_U101 ( .A(mult_50_n254), .B(mult_50_n252), .CI(mult_50_n261), 
        .CO(mult_50_n247), .S(mult_50_n248) );
  FA_X1 mult_50_U100 ( .A(mult_50_n259), .B(mult_50_n250), .CI(mult_50_n248), 
        .CO(mult_50_n245), .S(mult_50_n246) );
  FA_X1 mult_50_U97 ( .A(mult_50_n395), .B(mult_50_n359), .CI(mult_50_n408), 
        .CO(mult_50_n241), .S(mult_50_n242) );
  FA_X1 mult_50_U96 ( .A(mult_50_n335), .B(mult_50_n371), .CI(mult_50_n255), 
        .CO(mult_50_n239), .S(mult_50_n240) );
  FA_X1 mult_50_U95 ( .A(mult_50_n253), .B(mult_50_n244), .CI(mult_50_n251), 
        .CO(mult_50_n237), .S(mult_50_n238) );
  FA_X1 mult_50_U94 ( .A(mult_50_n240), .B(mult_50_n242), .CI(mult_50_n249), 
        .CO(mult_50_n235), .S(mult_50_n236) );
  FA_X1 mult_50_U93 ( .A(mult_50_n247), .B(mult_50_n238), .CI(mult_50_n236), 
        .CO(mult_50_n233), .S(mult_50_n234) );
  FA_X1 mult_50_U91 ( .A(mult_50_n382), .B(mult_50_n346), .CI(mult_50_n232), 
        .CO(mult_50_n229), .S(mult_50_n230) );
  FA_X1 mult_50_U90 ( .A(mult_50_n334), .B(mult_50_n370), .CI(mult_50_n358), 
        .CO(mult_50_n227), .S(mult_50_n228) );
  FA_X1 mult_50_U89 ( .A(mult_50_n241), .B(mult_50_n243), .CI(mult_50_n239), 
        .CO(mult_50_n225), .S(mult_50_n226) );
  FA_X1 mult_50_U88 ( .A(mult_50_n230), .B(mult_50_n228), .CI(mult_50_n237), 
        .CO(mult_50_n223), .S(mult_50_n224) );
  FA_X1 mult_50_U87 ( .A(mult_50_n235), .B(mult_50_n226), .CI(mult_50_n224), 
        .CO(mult_50_n221), .S(mult_50_n222) );
  FA_X1 mult_50_U86 ( .A(mult_50_n231), .B(mult_50_n333), .CI(mult_50_n394), 
        .CO(mult_50_n219), .S(mult_50_n220) );
  FA_X1 mult_50_U85 ( .A(mult_50_n345), .B(mult_50_n381), .CI(mult_50_n357), 
        .CO(mult_50_n217), .S(mult_50_n218) );
  FA_X1 mult_50_U84 ( .A(mult_50_n229), .B(mult_50_n369), .CI(mult_50_n227), 
        .CO(mult_50_n215), .S(mult_50_n216) );
  FA_X1 mult_50_U83 ( .A(mult_50_n220), .B(mult_50_n218), .CI(mult_50_n225), 
        .CO(mult_50_n213), .S(mult_50_n214) );
  FA_X1 mult_50_U82 ( .A(mult_50_n223), .B(mult_50_n216), .CI(mult_50_n214), 
        .CO(mult_50_n211), .S(mult_50_n212) );
  FA_X1 mult_50_U80 ( .A(mult_50_n368), .B(mult_50_n344), .CI(mult_50_n210), 
        .CO(mult_50_n207), .S(mult_50_n208) );
  FA_X1 mult_50_U79 ( .A(mult_50_n332), .B(mult_50_n356), .CI(mult_50_n219), 
        .CO(mult_50_n205), .S(mult_50_n206) );
  FA_X1 mult_50_U78 ( .A(mult_50_n208), .B(mult_50_n217), .CI(mult_50_n215), 
        .CO(mult_50_n203), .S(mult_50_n204) );
  FA_X1 mult_50_U77 ( .A(mult_50_n213), .B(mult_50_n206), .CI(mult_50_n204), 
        .CO(mult_50_n201), .S(mult_50_n202) );
  FA_X1 mult_50_U76 ( .A(mult_50_n209), .B(mult_50_n331), .CI(mult_50_n380), 
        .CO(mult_50_n199), .S(mult_50_n200) );
  FA_X1 mult_50_U75 ( .A(mult_50_n355), .B(mult_50_n343), .CI(mult_50_n367), 
        .CO(mult_50_n197), .S(mult_50_n198) );
  FA_X1 mult_50_U74 ( .A(mult_50_n198), .B(mult_50_n207), .CI(mult_50_n200), 
        .CO(mult_50_n195), .S(mult_50_n196) );
  FA_X1 mult_50_U73 ( .A(mult_50_n203), .B(mult_50_n205), .CI(mult_50_n196), 
        .CO(mult_50_n193), .S(mult_50_n194) );
  FA_X1 mult_50_U71 ( .A(mult_50_n330), .B(mult_50_n342), .CI(mult_50_n192), 
        .CO(mult_50_n189), .S(mult_50_n190) );
  FA_X1 mult_50_U70 ( .A(mult_50_n199), .B(mult_50_n354), .CI(mult_50_n197), 
        .CO(mult_50_n187), .S(mult_50_n188) );
  FA_X1 mult_50_U69 ( .A(mult_50_n188), .B(mult_50_n190), .CI(mult_50_n195), 
        .CO(mult_50_n185), .S(mult_50_n186) );
  FA_X1 mult_50_U68 ( .A(mult_50_n191), .B(mult_50_n329), .CI(mult_50_n366), 
        .CO(mult_50_n183), .S(mult_50_n184) );
  FA_X1 mult_50_U67 ( .A(mult_50_n341), .B(mult_50_n353), .CI(mult_50_n189), 
        .CO(mult_50_n181), .S(mult_50_n182) );
  FA_X1 mult_50_U66 ( .A(mult_50_n187), .B(mult_50_n184), .CI(mult_50_n182), 
        .CO(mult_50_n179), .S(mult_50_n180) );
  FA_X1 mult_50_U64 ( .A(mult_50_n328), .B(mult_50_n340), .CI(mult_50_n178), 
        .CO(mult_50_n175), .S(mult_50_n176) );
  FA_X1 mult_50_U63 ( .A(mult_50_n176), .B(mult_50_n183), .CI(mult_50_n181), 
        .CO(mult_50_n173), .S(mult_50_n174) );
  FA_X1 mult_50_U62 ( .A(mult_50_n327), .B(mult_50_n177), .CI(mult_50_n352), 
        .CO(mult_50_n171), .S(mult_50_n172) );
  FA_X1 mult_50_U61 ( .A(mult_50_n175), .B(mult_50_n339), .CI(mult_50_n172), 
        .CO(mult_50_n169), .S(mult_50_n170) );
  FA_X1 mult_50_U59 ( .A(mult_50_n168), .B(mult_50_n326), .CI(mult_50_n171), 
        .CO(mult_50_n165), .S(mult_50_n166) );
  FA_X1 mult_50_U58 ( .A(mult_50_n325), .B(mult_50_n167), .CI(mult_50_n338), 
        .CO(mult_50_n163), .S(mult_50_n164) );
  FA_X1 mult_50_U44 ( .A(mult_50_n246), .B(mult_50_n257), .CI(mult_50_n149), 
        .CO(mult_50_n148), .S(temp3_13_) );
  FA_X1 mult_50_U43 ( .A(mult_50_n234), .B(mult_50_n245), .CI(mult_50_n148), 
        .CO(mult_50_n147), .S(temp3_14_) );
  FA_X1 mult_50_U42 ( .A(mult_50_n222), .B(mult_50_n233), .CI(mult_50_n147), 
        .CO(mult_50_n146), .S(temp3_15_) );
  FA_X1 mult_50_U41 ( .A(mult_50_n212), .B(mult_50_n221), .CI(mult_50_n146), 
        .CO(mult_50_n145), .S(temp3_16_) );
  FA_X1 mult_50_U40 ( .A(mult_50_n202), .B(mult_50_n211), .CI(mult_50_n145), 
        .CO(mult_50_n144), .S(temp3_17_) );
  FA_X1 mult_50_U39 ( .A(mult_50_n194), .B(mult_50_n201), .CI(mult_50_n144), 
        .CO(mult_50_n143), .S(temp3_18_) );
  FA_X1 mult_50_U38 ( .A(mult_50_n186), .B(mult_50_n193), .CI(mult_50_n143), 
        .CO(mult_50_n142), .S(temp3_19_) );
  FA_X1 mult_50_U37 ( .A(mult_50_n180), .B(mult_50_n185), .CI(mult_50_n142), 
        .CO(mult_50_n141), .S(temp3_20_) );
  FA_X1 mult_50_U30 ( .A(mult_50_n174), .B(mult_50_n179), .CI(mult_50_n141), 
        .CO(mult_50_n140), .S(temp3_21_) );
  FA_X1 mult_50_U20 ( .A(mult_50_n170), .B(mult_50_n173), .CI(mult_50_n140), 
        .CO(mult_50_n139), .S(temp3_22_) );
  FA_X1 mult_50_U10 ( .A(mult_50_n166), .B(mult_50_n169), .CI(mult_50_n139), 
        .CO(mult_50_n138), .S(temp3_23_) );
  FA_X1 mult_50_U9 ( .A(mult_50_n165), .B(mult_50_n164), .CI(mult_50_n138), 
        .CO(mult_50_n137), .S(temp3_24_) );
  FA_X1 mult_50_U8 ( .A(mult_50_n163), .B(mult_50_n162), .CI(mult_50_n137), 
        .CO(mult_50_n136), .S(temp3_25_) );
  XOR2_X1 mult_52_U691 ( .A(reg2[2]), .B(n158), .Z(mult_52_n798) );
  NOR2_X1 mult_52_U690 ( .A1(mult_52_n635), .A2(B2[1]), .ZN(mult_52_n803) );
  INV_X1 mult_52_U689 ( .A(mult_52_n803), .ZN(mult_52_n805) );
  NAND2_X1 mult_52_U688 ( .A1(n158), .A2(mult_52_n650), .ZN(mult_52_n648) );
  XNOR2_X1 mult_52_U687 ( .A(B2[2]), .B(n158), .ZN(mult_52_n647) );
  OAI22_X1 mult_52_U686 ( .A1(mult_52_n805), .A2(mult_52_n648), .B1(
        mult_52_n647), .B2(mult_52_n650), .ZN(mult_52_n804) );
  NAND2_X1 mult_52_U685 ( .A1(mult_52_n798), .A2(mult_52_n804), .ZN(
        mult_52_n801) );
  NAND2_X1 mult_52_U684 ( .A1(mult_52_n803), .A2(mult_52_n804), .ZN(
        mult_52_n802) );
  INV_X1 mult_52_U683 ( .A(B2[0]), .ZN(mult_52_n679) );
  MUX2_X1 mult_52_U682 ( .A(mult_52_n801), .B(mult_52_n802), .S(mult_52_n679), 
        .Z(mult_52_n800) );
  INV_X1 mult_52_U681 ( .A(mult_52_n800), .ZN(mult_52_n795) );
  XNOR2_X1 mult_52_U680 ( .A(mult_52_n636), .B(reg2[2]), .ZN(mult_52_n799) );
  NAND2_X1 mult_52_U679 ( .A1(mult_52_n664), .A2(mult_52_n799), .ZN(
        mult_52_n663) );
  NAND3_X1 mult_52_U678 ( .A1(mult_52_n798), .A2(mult_52_n679), .A3(n160), 
        .ZN(mult_52_n797) );
  OAI21_X1 mult_52_U677 ( .B1(mult_52_n636), .B2(mult_52_n663), .A(
        mult_52_n797), .ZN(mult_52_n796) );
  AOI222_X1 mult_52_U676 ( .A1(mult_52_n795), .A2(mult_52_n316), .B1(
        mult_52_n796), .B2(mult_52_n795), .C1(mult_52_n796), .C2(mult_52_n316), 
        .ZN(mult_52_n794) );
  INV_X1 mult_52_U675 ( .A(mult_52_n794), .ZN(mult_52_n793) );
  AOI222_X1 mult_52_U674 ( .A1(mult_52_n793), .A2(mult_52_n314), .B1(
        mult_52_n793), .B2(mult_52_n315), .C1(mult_52_n315), .C2(mult_52_n314), 
        .ZN(mult_52_n792) );
  INV_X1 mult_52_U673 ( .A(mult_52_n792), .ZN(mult_52_n791) );
  AOI222_X1 mult_52_U672 ( .A1(mult_52_n791), .A2(mult_52_n310), .B1(
        mult_52_n791), .B2(mult_52_n313), .C1(mult_52_n313), .C2(mult_52_n310), 
        .ZN(mult_52_n790) );
  INV_X1 mult_52_U671 ( .A(mult_52_n790), .ZN(mult_52_n789) );
  AOI222_X1 mult_52_U670 ( .A1(mult_52_n789), .A2(mult_52_n306), .B1(
        mult_52_n789), .B2(mult_52_n309), .C1(mult_52_n309), .C2(mult_52_n306), 
        .ZN(mult_52_n788) );
  INV_X1 mult_52_U669 ( .A(mult_52_n788), .ZN(mult_52_n787) );
  AOI222_X1 mult_52_U668 ( .A1(mult_52_n787), .A2(mult_52_n300), .B1(
        mult_52_n787), .B2(mult_52_n305), .C1(mult_52_n305), .C2(mult_52_n300), 
        .ZN(mult_52_n786) );
  INV_X1 mult_52_U667 ( .A(mult_52_n786), .ZN(mult_52_n785) );
  AOI222_X1 mult_52_U666 ( .A1(mult_52_n785), .A2(mult_52_n294), .B1(
        mult_52_n785), .B2(mult_52_n299), .C1(mult_52_n299), .C2(mult_52_n294), 
        .ZN(mult_52_n784) );
  INV_X1 mult_52_U665 ( .A(mult_52_n784), .ZN(mult_52_n783) );
  AOI222_X1 mult_52_U664 ( .A1(mult_52_n783), .A2(mult_52_n286), .B1(
        mult_52_n783), .B2(mult_52_n293), .C1(mult_52_n293), .C2(mult_52_n286), 
        .ZN(mult_52_n780) );
  INV_X1 mult_52_U663 ( .A(mult_52_n278), .ZN(mult_52_n781) );
  INV_X1 mult_52_U662 ( .A(mult_52_n285), .ZN(mult_52_n782) );
  OAI222_X1 mult_52_U661 ( .A1(mult_52_n780), .A2(mult_52_n781), .B1(
        mult_52_n780), .B2(mult_52_n782), .C1(mult_52_n782), .C2(mult_52_n781), 
        .ZN(mult_52_n779) );
  AOI222_X1 mult_52_U660 ( .A1(mult_52_n779), .A2(mult_52_n268), .B1(
        mult_52_n779), .B2(mult_52_n277), .C1(mult_52_n277), .C2(mult_52_n268), 
        .ZN(mult_52_n776) );
  INV_X1 mult_52_U659 ( .A(mult_52_n258), .ZN(mult_52_n777) );
  INV_X1 mult_52_U658 ( .A(mult_52_n267), .ZN(mult_52_n778) );
  OAI222_X1 mult_52_U657 ( .A1(mult_52_n776), .A2(mult_52_n777), .B1(
        mult_52_n776), .B2(mult_52_n778), .C1(mult_52_n778), .C2(mult_52_n777), 
        .ZN(mult_52_n149) );
  XOR2_X1 mult_52_U656 ( .A(B2[12]), .B(n170), .Z(mult_52_n763) );
  XNOR2_X1 mult_52_U655 ( .A(mult_52_n641), .B(reg2[12]), .ZN(mult_52_n775) );
  NAND2_X1 mult_52_U654 ( .A1(mult_52_n748), .A2(mult_52_n775), .ZN(
        mult_52_n750) );
  INV_X1 mult_52_U653 ( .A(mult_52_n750), .ZN(mult_52_n644) );
  INV_X1 mult_52_U652 ( .A(mult_52_n748), .ZN(mult_52_n645) );
  XNOR2_X1 mult_52_U651 ( .A(B2[13]), .B(mult_52_n641), .ZN(mult_52_n646) );
  AOI22_X1 mult_52_U650 ( .A1(mult_52_n763), .A2(mult_52_n644), .B1(
        mult_52_n645), .B2(mult_52_n646), .ZN(mult_52_n162) );
  XNOR2_X1 mult_52_U649 ( .A(B2[12]), .B(n168), .ZN(mult_52_n745) );
  XNOR2_X1 mult_52_U648 ( .A(mult_52_n640), .B(reg2[10]), .ZN(mult_52_n774) );
  NAND2_X1 mult_52_U647 ( .A1(mult_52_n731), .A2(mult_52_n774), .ZN(
        mult_52_n733) );
  XNOR2_X1 mult_52_U646 ( .A(B2[13]), .B(n168), .ZN(mult_52_n747) );
  OAI22_X1 mult_52_U645 ( .A1(mult_52_n745), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n747), .ZN(mult_52_n167) );
  INV_X1 mult_52_U644 ( .A(mult_52_n167), .ZN(mult_52_n168) );
  XNOR2_X1 mult_52_U643 ( .A(B2[12]), .B(n166), .ZN(mult_52_n728) );
  XNOR2_X1 mult_52_U642 ( .A(mult_52_n639), .B(reg2[8]), .ZN(mult_52_n773) );
  NAND2_X1 mult_52_U641 ( .A1(mult_52_n714), .A2(mult_52_n773), .ZN(
        mult_52_n716) );
  XNOR2_X1 mult_52_U640 ( .A(B2[13]), .B(n166), .ZN(mult_52_n730) );
  OAI22_X1 mult_52_U639 ( .A1(mult_52_n728), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n730), .ZN(mult_52_n177) );
  INV_X1 mult_52_U638 ( .A(mult_52_n177), .ZN(mult_52_n178) );
  XNOR2_X1 mult_52_U637 ( .A(B2[12]), .B(n164), .ZN(mult_52_n711) );
  XNOR2_X1 mult_52_U636 ( .A(mult_52_n638), .B(reg2[6]), .ZN(mult_52_n772) );
  NAND2_X1 mult_52_U635 ( .A1(mult_52_n697), .A2(mult_52_n772), .ZN(
        mult_52_n699) );
  XNOR2_X1 mult_52_U634 ( .A(B2[13]), .B(n164), .ZN(mult_52_n713) );
  OAI22_X1 mult_52_U633 ( .A1(mult_52_n711), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n713), .ZN(mult_52_n191) );
  INV_X1 mult_52_U632 ( .A(mult_52_n191), .ZN(mult_52_n192) );
  XNOR2_X1 mult_52_U631 ( .A(B2[12]), .B(n162), .ZN(mult_52_n694) );
  XNOR2_X1 mult_52_U630 ( .A(mult_52_n637), .B(reg2[4]), .ZN(mult_52_n771) );
  NAND2_X1 mult_52_U629 ( .A1(mult_52_n680), .A2(mult_52_n771), .ZN(
        mult_52_n682) );
  XNOR2_X1 mult_52_U628 ( .A(B2[13]), .B(n162), .ZN(mult_52_n696) );
  OAI22_X1 mult_52_U627 ( .A1(mult_52_n694), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n696), .ZN(mult_52_n209) );
  INV_X1 mult_52_U626 ( .A(mult_52_n209), .ZN(mult_52_n210) );
  XNOR2_X1 mult_52_U625 ( .A(B2[12]), .B(n160), .ZN(mult_52_n676) );
  XNOR2_X1 mult_52_U624 ( .A(B2[13]), .B(n160), .ZN(mult_52_n678) );
  OAI22_X1 mult_52_U623 ( .A1(mult_52_n676), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n678), .ZN(mult_52_n231) );
  INV_X1 mult_52_U622 ( .A(mult_52_n231), .ZN(mult_52_n232) );
  XNOR2_X1 mult_52_U621 ( .A(B2[3]), .B(n168), .ZN(mult_52_n736) );
  XNOR2_X1 mult_52_U620 ( .A(B2[4]), .B(n168), .ZN(mult_52_n737) );
  OAI22_X1 mult_52_U619 ( .A1(mult_52_n736), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n737), .ZN(mult_52_n769) );
  XNOR2_X1 mult_52_U618 ( .A(B2[9]), .B(n162), .ZN(mult_52_n691) );
  XNOR2_X1 mult_52_U617 ( .A(B2[10]), .B(n162), .ZN(mult_52_n692) );
  OAI22_X1 mult_52_U616 ( .A1(mult_52_n691), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n692), .ZN(mult_52_n770) );
  OR2_X1 mult_52_U615 ( .A1(mult_52_n769), .A2(mult_52_n770), .ZN(mult_52_n243) );
  XNOR2_X1 mult_52_U614 ( .A(mult_52_n769), .B(mult_52_n770), .ZN(mult_52_n244) );
  NAND3_X1 mult_52_U613 ( .A1(mult_52_n645), .A2(mult_52_n679), .A3(n170), 
        .ZN(mult_52_n768) );
  OAI21_X1 mult_52_U612 ( .B1(mult_52_n641), .B2(mult_52_n750), .A(
        mult_52_n768), .ZN(mult_52_n317) );
  OR3_X1 mult_52_U611 ( .A1(mult_52_n731), .A2(B2[0]), .A3(mult_52_n640), .ZN(
        mult_52_n767) );
  OAI21_X1 mult_52_U610 ( .B1(mult_52_n640), .B2(mult_52_n733), .A(
        mult_52_n767), .ZN(mult_52_n318) );
  OR3_X1 mult_52_U609 ( .A1(mult_52_n714), .A2(B2[0]), .A3(mult_52_n639), .ZN(
        mult_52_n766) );
  OAI21_X1 mult_52_U608 ( .B1(mult_52_n639), .B2(mult_52_n716), .A(
        mult_52_n766), .ZN(mult_52_n319) );
  OR3_X1 mult_52_U607 ( .A1(mult_52_n697), .A2(B2[0]), .A3(mult_52_n638), .ZN(
        mult_52_n765) );
  OAI21_X1 mult_52_U606 ( .B1(mult_52_n638), .B2(mult_52_n699), .A(
        mult_52_n765), .ZN(mult_52_n320) );
  OR3_X1 mult_52_U605 ( .A1(mult_52_n680), .A2(B2[0]), .A3(mult_52_n637), .ZN(
        mult_52_n764) );
  OAI21_X1 mult_52_U604 ( .B1(mult_52_n637), .B2(mult_52_n682), .A(
        mult_52_n764), .ZN(mult_52_n321) );
  XNOR2_X1 mult_52_U603 ( .A(B2[11]), .B(n170), .ZN(mult_52_n761) );
  INV_X1 mult_52_U602 ( .A(mult_52_n763), .ZN(mult_52_n762) );
  OAI22_X1 mult_52_U601 ( .A1(mult_52_n761), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n762), .ZN(mult_52_n325) );
  XNOR2_X1 mult_52_U600 ( .A(B2[10]), .B(n170), .ZN(mult_52_n760) );
  OAI22_X1 mult_52_U599 ( .A1(mult_52_n760), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n761), .ZN(mult_52_n326) );
  XNOR2_X1 mult_52_U598 ( .A(B2[9]), .B(n170), .ZN(mult_52_n759) );
  OAI22_X1 mult_52_U597 ( .A1(mult_52_n759), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n760), .ZN(mult_52_n327) );
  XNOR2_X1 mult_52_U596 ( .A(B2[8]), .B(n170), .ZN(mult_52_n758) );
  OAI22_X1 mult_52_U595 ( .A1(mult_52_n758), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n759), .ZN(mult_52_n328) );
  XNOR2_X1 mult_52_U594 ( .A(B2[7]), .B(n170), .ZN(mult_52_n757) );
  OAI22_X1 mult_52_U593 ( .A1(mult_52_n757), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n758), .ZN(mult_52_n329) );
  XNOR2_X1 mult_52_U592 ( .A(B2[6]), .B(n170), .ZN(mult_52_n756) );
  OAI22_X1 mult_52_U591 ( .A1(mult_52_n756), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n757), .ZN(mult_52_n330) );
  XNOR2_X1 mult_52_U590 ( .A(B2[5]), .B(n170), .ZN(mult_52_n755) );
  OAI22_X1 mult_52_U589 ( .A1(mult_52_n755), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n756), .ZN(mult_52_n331) );
  XNOR2_X1 mult_52_U588 ( .A(B2[4]), .B(n170), .ZN(mult_52_n754) );
  OAI22_X1 mult_52_U587 ( .A1(mult_52_n754), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n755), .ZN(mult_52_n332) );
  XNOR2_X1 mult_52_U586 ( .A(B2[3]), .B(n170), .ZN(mult_52_n753) );
  OAI22_X1 mult_52_U585 ( .A1(mult_52_n753), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n754), .ZN(mult_52_n333) );
  XNOR2_X1 mult_52_U584 ( .A(B2[2]), .B(n170), .ZN(mult_52_n752) );
  OAI22_X1 mult_52_U583 ( .A1(mult_52_n752), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n753), .ZN(mult_52_n334) );
  XNOR2_X1 mult_52_U582 ( .A(B2[1]), .B(n170), .ZN(mult_52_n751) );
  OAI22_X1 mult_52_U581 ( .A1(mult_52_n751), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n752), .ZN(mult_52_n335) );
  XNOR2_X1 mult_52_U580 ( .A(n170), .B(B2[0]), .ZN(mult_52_n749) );
  OAI22_X1 mult_52_U579 ( .A1(mult_52_n749), .A2(mult_52_n750), .B1(
        mult_52_n748), .B2(mult_52_n751), .ZN(mult_52_n336) );
  NOR2_X1 mult_52_U578 ( .A1(mult_52_n679), .A2(mult_52_n748), .ZN(
        mult_52_n337) );
  AOI21_X1 mult_52_U577 ( .B1(mult_52_n733), .B2(mult_52_n731), .A(
        mult_52_n747), .ZN(mult_52_n746) );
  INV_X1 mult_52_U576 ( .A(mult_52_n746), .ZN(mult_52_n338) );
  XNOR2_X1 mult_52_U575 ( .A(B2[11]), .B(n168), .ZN(mult_52_n744) );
  OAI22_X1 mult_52_U574 ( .A1(mult_52_n744), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n745), .ZN(mult_52_n339) );
  XNOR2_X1 mult_52_U573 ( .A(B2[10]), .B(n168), .ZN(mult_52_n743) );
  OAI22_X1 mult_52_U572 ( .A1(mult_52_n743), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n744), .ZN(mult_52_n340) );
  XNOR2_X1 mult_52_U571 ( .A(B2[9]), .B(n168), .ZN(mult_52_n742) );
  OAI22_X1 mult_52_U570 ( .A1(mult_52_n742), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n743), .ZN(mult_52_n341) );
  XNOR2_X1 mult_52_U569 ( .A(B2[8]), .B(n168), .ZN(mult_52_n741) );
  OAI22_X1 mult_52_U568 ( .A1(mult_52_n741), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n742), .ZN(mult_52_n342) );
  XNOR2_X1 mult_52_U567 ( .A(B2[7]), .B(n168), .ZN(mult_52_n740) );
  OAI22_X1 mult_52_U566 ( .A1(mult_52_n740), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n741), .ZN(mult_52_n343) );
  XNOR2_X1 mult_52_U565 ( .A(B2[6]), .B(n168), .ZN(mult_52_n739) );
  OAI22_X1 mult_52_U564 ( .A1(mult_52_n739), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n740), .ZN(mult_52_n344) );
  XNOR2_X1 mult_52_U563 ( .A(B2[5]), .B(n168), .ZN(mult_52_n738) );
  OAI22_X1 mult_52_U562 ( .A1(mult_52_n738), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n739), .ZN(mult_52_n345) );
  OAI22_X1 mult_52_U561 ( .A1(mult_52_n737), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n738), .ZN(mult_52_n346) );
  XNOR2_X1 mult_52_U560 ( .A(B2[2]), .B(n168), .ZN(mult_52_n735) );
  OAI22_X1 mult_52_U559 ( .A1(mult_52_n735), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n736), .ZN(mult_52_n348) );
  XNOR2_X1 mult_52_U558 ( .A(B2[1]), .B(n168), .ZN(mult_52_n734) );
  OAI22_X1 mult_52_U557 ( .A1(mult_52_n734), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n735), .ZN(mult_52_n349) );
  XNOR2_X1 mult_52_U556 ( .A(n168), .B(B2[0]), .ZN(mult_52_n732) );
  OAI22_X1 mult_52_U555 ( .A1(mult_52_n732), .A2(mult_52_n733), .B1(
        mult_52_n731), .B2(mult_52_n734), .ZN(mult_52_n350) );
  NOR2_X1 mult_52_U554 ( .A1(mult_52_n679), .A2(mult_52_n731), .ZN(
        mult_52_n351) );
  AOI21_X1 mult_52_U553 ( .B1(mult_52_n716), .B2(mult_52_n714), .A(
        mult_52_n730), .ZN(mult_52_n729) );
  INV_X1 mult_52_U552 ( .A(mult_52_n729), .ZN(mult_52_n352) );
  XNOR2_X1 mult_52_U551 ( .A(B2[11]), .B(n166), .ZN(mult_52_n727) );
  OAI22_X1 mult_52_U550 ( .A1(mult_52_n727), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n728), .ZN(mult_52_n353) );
  XNOR2_X1 mult_52_U549 ( .A(B2[10]), .B(n166), .ZN(mult_52_n726) );
  OAI22_X1 mult_52_U548 ( .A1(mult_52_n726), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n727), .ZN(mult_52_n354) );
  XNOR2_X1 mult_52_U547 ( .A(B2[9]), .B(n166), .ZN(mult_52_n725) );
  OAI22_X1 mult_52_U546 ( .A1(mult_52_n725), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n726), .ZN(mult_52_n355) );
  XNOR2_X1 mult_52_U545 ( .A(B2[8]), .B(n166), .ZN(mult_52_n724) );
  OAI22_X1 mult_52_U544 ( .A1(mult_52_n724), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n725), .ZN(mult_52_n356) );
  XNOR2_X1 mult_52_U543 ( .A(B2[7]), .B(n166), .ZN(mult_52_n723) );
  OAI22_X1 mult_52_U542 ( .A1(mult_52_n723), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n724), .ZN(mult_52_n357) );
  XNOR2_X1 mult_52_U541 ( .A(B2[6]), .B(n166), .ZN(mult_52_n722) );
  OAI22_X1 mult_52_U540 ( .A1(mult_52_n722), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n723), .ZN(mult_52_n358) );
  XNOR2_X1 mult_52_U539 ( .A(B2[5]), .B(n166), .ZN(mult_52_n721) );
  OAI22_X1 mult_52_U538 ( .A1(mult_52_n721), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n722), .ZN(mult_52_n359) );
  XNOR2_X1 mult_52_U537 ( .A(B2[4]), .B(n166), .ZN(mult_52_n720) );
  OAI22_X1 mult_52_U536 ( .A1(mult_52_n720), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n721), .ZN(mult_52_n360) );
  XNOR2_X1 mult_52_U535 ( .A(B2[3]), .B(n166), .ZN(mult_52_n719) );
  OAI22_X1 mult_52_U534 ( .A1(mult_52_n719), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n720), .ZN(mult_52_n361) );
  XNOR2_X1 mult_52_U533 ( .A(B2[2]), .B(n166), .ZN(mult_52_n718) );
  OAI22_X1 mult_52_U532 ( .A1(mult_52_n718), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n719), .ZN(mult_52_n362) );
  XNOR2_X1 mult_52_U531 ( .A(B2[1]), .B(n166), .ZN(mult_52_n717) );
  OAI22_X1 mult_52_U530 ( .A1(mult_52_n717), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n718), .ZN(mult_52_n363) );
  XNOR2_X1 mult_52_U529 ( .A(n166), .B(B2[0]), .ZN(mult_52_n715) );
  OAI22_X1 mult_52_U528 ( .A1(mult_52_n715), .A2(mult_52_n716), .B1(
        mult_52_n714), .B2(mult_52_n717), .ZN(mult_52_n364) );
  NOR2_X1 mult_52_U527 ( .A1(mult_52_n679), .A2(mult_52_n714), .ZN(
        mult_52_n365) );
  AOI21_X1 mult_52_U526 ( .B1(mult_52_n699), .B2(mult_52_n697), .A(
        mult_52_n713), .ZN(mult_52_n712) );
  INV_X1 mult_52_U525 ( .A(mult_52_n712), .ZN(mult_52_n366) );
  XNOR2_X1 mult_52_U524 ( .A(B2[11]), .B(n164), .ZN(mult_52_n710) );
  OAI22_X1 mult_52_U523 ( .A1(mult_52_n710), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n711), .ZN(mult_52_n367) );
  XNOR2_X1 mult_52_U522 ( .A(B2[10]), .B(n164), .ZN(mult_52_n709) );
  OAI22_X1 mult_52_U521 ( .A1(mult_52_n709), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n710), .ZN(mult_52_n368) );
  XNOR2_X1 mult_52_U520 ( .A(B2[9]), .B(n164), .ZN(mult_52_n708) );
  OAI22_X1 mult_52_U519 ( .A1(mult_52_n708), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n709), .ZN(mult_52_n369) );
  XNOR2_X1 mult_52_U518 ( .A(B2[8]), .B(n164), .ZN(mult_52_n707) );
  OAI22_X1 mult_52_U517 ( .A1(mult_52_n707), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n708), .ZN(mult_52_n370) );
  XNOR2_X1 mult_52_U516 ( .A(B2[7]), .B(n164), .ZN(mult_52_n706) );
  OAI22_X1 mult_52_U515 ( .A1(mult_52_n706), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n707), .ZN(mult_52_n371) );
  XNOR2_X1 mult_52_U514 ( .A(B2[6]), .B(n164), .ZN(mult_52_n705) );
  OAI22_X1 mult_52_U513 ( .A1(mult_52_n705), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n706), .ZN(mult_52_n372) );
  XNOR2_X1 mult_52_U512 ( .A(B2[5]), .B(n164), .ZN(mult_52_n704) );
  OAI22_X1 mult_52_U511 ( .A1(mult_52_n704), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n705), .ZN(mult_52_n373) );
  XNOR2_X1 mult_52_U510 ( .A(B2[4]), .B(n164), .ZN(mult_52_n703) );
  OAI22_X1 mult_52_U509 ( .A1(mult_52_n703), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n704), .ZN(mult_52_n374) );
  XNOR2_X1 mult_52_U508 ( .A(B2[3]), .B(n164), .ZN(mult_52_n702) );
  OAI22_X1 mult_52_U507 ( .A1(mult_52_n702), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n703), .ZN(mult_52_n375) );
  XNOR2_X1 mult_52_U506 ( .A(B2[2]), .B(n164), .ZN(mult_52_n701) );
  OAI22_X1 mult_52_U505 ( .A1(mult_52_n701), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n702), .ZN(mult_52_n376) );
  XNOR2_X1 mult_52_U504 ( .A(B2[1]), .B(n164), .ZN(mult_52_n700) );
  OAI22_X1 mult_52_U503 ( .A1(mult_52_n700), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n701), .ZN(mult_52_n377) );
  XNOR2_X1 mult_52_U502 ( .A(n164), .B(B2[0]), .ZN(mult_52_n698) );
  OAI22_X1 mult_52_U501 ( .A1(mult_52_n698), .A2(mult_52_n699), .B1(
        mult_52_n697), .B2(mult_52_n700), .ZN(mult_52_n378) );
  NOR2_X1 mult_52_U500 ( .A1(mult_52_n679), .A2(mult_52_n697), .ZN(
        mult_52_n379) );
  AOI21_X1 mult_52_U499 ( .B1(mult_52_n682), .B2(mult_52_n680), .A(
        mult_52_n696), .ZN(mult_52_n695) );
  INV_X1 mult_52_U498 ( .A(mult_52_n695), .ZN(mult_52_n380) );
  XNOR2_X1 mult_52_U497 ( .A(B2[11]), .B(n162), .ZN(mult_52_n693) );
  OAI22_X1 mult_52_U496 ( .A1(mult_52_n693), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n694), .ZN(mult_52_n381) );
  OAI22_X1 mult_52_U495 ( .A1(mult_52_n692), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n693), .ZN(mult_52_n382) );
  XNOR2_X1 mult_52_U494 ( .A(B2[8]), .B(n162), .ZN(mult_52_n690) );
  OAI22_X1 mult_52_U493 ( .A1(mult_52_n690), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n691), .ZN(mult_52_n384) );
  XNOR2_X1 mult_52_U492 ( .A(B2[7]), .B(n162), .ZN(mult_52_n689) );
  OAI22_X1 mult_52_U491 ( .A1(mult_52_n689), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n690), .ZN(mult_52_n385) );
  XNOR2_X1 mult_52_U490 ( .A(B2[6]), .B(n162), .ZN(mult_52_n688) );
  OAI22_X1 mult_52_U489 ( .A1(mult_52_n688), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n689), .ZN(mult_52_n386) );
  XNOR2_X1 mult_52_U488 ( .A(B2[5]), .B(n162), .ZN(mult_52_n687) );
  OAI22_X1 mult_52_U487 ( .A1(mult_52_n687), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n688), .ZN(mult_52_n387) );
  XNOR2_X1 mult_52_U486 ( .A(B2[4]), .B(n162), .ZN(mult_52_n686) );
  OAI22_X1 mult_52_U485 ( .A1(mult_52_n686), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n687), .ZN(mult_52_n388) );
  XNOR2_X1 mult_52_U484 ( .A(B2[3]), .B(n162), .ZN(mult_52_n685) );
  OAI22_X1 mult_52_U483 ( .A1(mult_52_n685), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n686), .ZN(mult_52_n389) );
  XNOR2_X1 mult_52_U482 ( .A(B2[2]), .B(n162), .ZN(mult_52_n684) );
  OAI22_X1 mult_52_U481 ( .A1(mult_52_n684), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n685), .ZN(mult_52_n390) );
  XNOR2_X1 mult_52_U480 ( .A(B2[1]), .B(n162), .ZN(mult_52_n683) );
  OAI22_X1 mult_52_U479 ( .A1(mult_52_n683), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n684), .ZN(mult_52_n391) );
  XNOR2_X1 mult_52_U478 ( .A(n162), .B(B2[0]), .ZN(mult_52_n681) );
  OAI22_X1 mult_52_U477 ( .A1(mult_52_n681), .A2(mult_52_n682), .B1(
        mult_52_n680), .B2(mult_52_n683), .ZN(mult_52_n392) );
  NOR2_X1 mult_52_U476 ( .A1(mult_52_n679), .A2(mult_52_n680), .ZN(
        mult_52_n393) );
  AOI21_X1 mult_52_U475 ( .B1(mult_52_n663), .B2(mult_52_n664), .A(
        mult_52_n678), .ZN(mult_52_n677) );
  INV_X1 mult_52_U474 ( .A(mult_52_n677), .ZN(mult_52_n394) );
  XNOR2_X1 mult_52_U473 ( .A(B2[11]), .B(n160), .ZN(mult_52_n675) );
  OAI22_X1 mult_52_U472 ( .A1(mult_52_n675), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n676), .ZN(mult_52_n395) );
  XNOR2_X1 mult_52_U471 ( .A(B2[10]), .B(n160), .ZN(mult_52_n674) );
  OAI22_X1 mult_52_U470 ( .A1(mult_52_n674), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n675), .ZN(mult_52_n396) );
  XNOR2_X1 mult_52_U469 ( .A(B2[9]), .B(n160), .ZN(mult_52_n673) );
  OAI22_X1 mult_52_U468 ( .A1(mult_52_n673), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n674), .ZN(mult_52_n397) );
  XNOR2_X1 mult_52_U467 ( .A(B2[8]), .B(n160), .ZN(mult_52_n672) );
  OAI22_X1 mult_52_U466 ( .A1(mult_52_n672), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n673), .ZN(mult_52_n398) );
  XNOR2_X1 mult_52_U465 ( .A(B2[7]), .B(n160), .ZN(mult_52_n671) );
  OAI22_X1 mult_52_U464 ( .A1(mult_52_n671), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n672), .ZN(mult_52_n399) );
  XNOR2_X1 mult_52_U463 ( .A(B2[6]), .B(n160), .ZN(mult_52_n670) );
  OAI22_X1 mult_52_U462 ( .A1(mult_52_n670), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n671), .ZN(mult_52_n400) );
  XNOR2_X1 mult_52_U461 ( .A(B2[5]), .B(n160), .ZN(mult_52_n669) );
  OAI22_X1 mult_52_U460 ( .A1(mult_52_n669), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n670), .ZN(mult_52_n401) );
  XNOR2_X1 mult_52_U459 ( .A(B2[4]), .B(n160), .ZN(mult_52_n668) );
  OAI22_X1 mult_52_U458 ( .A1(mult_52_n668), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n669), .ZN(mult_52_n402) );
  XNOR2_X1 mult_52_U457 ( .A(B2[3]), .B(n160), .ZN(mult_52_n667) );
  OAI22_X1 mult_52_U456 ( .A1(mult_52_n667), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n668), .ZN(mult_52_n403) );
  XNOR2_X1 mult_52_U455 ( .A(B2[2]), .B(n160), .ZN(mult_52_n666) );
  OAI22_X1 mult_52_U454 ( .A1(mult_52_n666), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n667), .ZN(mult_52_n404) );
  XNOR2_X1 mult_52_U453 ( .A(B2[1]), .B(n160), .ZN(mult_52_n665) );
  OAI22_X1 mult_52_U452 ( .A1(mult_52_n665), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n666), .ZN(mult_52_n405) );
  XNOR2_X1 mult_52_U451 ( .A(n160), .B(B2[0]), .ZN(mult_52_n662) );
  OAI22_X1 mult_52_U450 ( .A1(mult_52_n662), .A2(mult_52_n663), .B1(
        mult_52_n664), .B2(mult_52_n665), .ZN(mult_52_n406) );
  XOR2_X1 mult_52_U449 ( .A(B2[13]), .B(mult_52_n635), .Z(mult_52_n660) );
  AOI21_X1 mult_52_U448 ( .B1(mult_52_n648), .B2(mult_52_n650), .A(
        mult_52_n660), .ZN(mult_52_n661) );
  INV_X1 mult_52_U447 ( .A(mult_52_n661), .ZN(mult_52_n408) );
  XNOR2_X1 mult_52_U446 ( .A(B2[12]), .B(n158), .ZN(mult_52_n659) );
  OAI22_X1 mult_52_U445 ( .A1(mult_52_n659), .A2(mult_52_n648), .B1(
        mult_52_n660), .B2(mult_52_n650), .ZN(mult_52_n409) );
  XNOR2_X1 mult_52_U444 ( .A(B2[11]), .B(n158), .ZN(mult_52_n658) );
  OAI22_X1 mult_52_U443 ( .A1(mult_52_n658), .A2(mult_52_n648), .B1(
        mult_52_n659), .B2(mult_52_n650), .ZN(mult_52_n410) );
  XNOR2_X1 mult_52_U442 ( .A(B2[10]), .B(n158), .ZN(mult_52_n657) );
  OAI22_X1 mult_52_U441 ( .A1(mult_52_n657), .A2(mult_52_n648), .B1(
        mult_52_n658), .B2(mult_52_n650), .ZN(mult_52_n411) );
  XNOR2_X1 mult_52_U440 ( .A(B2[9]), .B(n158), .ZN(mult_52_n656) );
  OAI22_X1 mult_52_U439 ( .A1(mult_52_n656), .A2(mult_52_n648), .B1(
        mult_52_n657), .B2(mult_52_n650), .ZN(mult_52_n412) );
  XNOR2_X1 mult_52_U438 ( .A(B2[8]), .B(n158), .ZN(mult_52_n655) );
  OAI22_X1 mult_52_U437 ( .A1(mult_52_n655), .A2(mult_52_n648), .B1(
        mult_52_n656), .B2(mult_52_n650), .ZN(mult_52_n413) );
  XNOR2_X1 mult_52_U436 ( .A(B2[7]), .B(n158), .ZN(mult_52_n654) );
  OAI22_X1 mult_52_U435 ( .A1(mult_52_n654), .A2(mult_52_n648), .B1(
        mult_52_n655), .B2(mult_52_n650), .ZN(mult_52_n414) );
  XNOR2_X1 mult_52_U434 ( .A(B2[6]), .B(n158), .ZN(mult_52_n653) );
  OAI22_X1 mult_52_U433 ( .A1(mult_52_n653), .A2(mult_52_n648), .B1(
        mult_52_n654), .B2(mult_52_n650), .ZN(mult_52_n415) );
  XNOR2_X1 mult_52_U432 ( .A(B2[5]), .B(n158), .ZN(mult_52_n652) );
  OAI22_X1 mult_52_U431 ( .A1(mult_52_n652), .A2(mult_52_n648), .B1(
        mult_52_n653), .B2(mult_52_n650), .ZN(mult_52_n416) );
  XNOR2_X1 mult_52_U430 ( .A(B2[4]), .B(n158), .ZN(mult_52_n651) );
  OAI22_X1 mult_52_U429 ( .A1(mult_52_n651), .A2(mult_52_n648), .B1(
        mult_52_n652), .B2(mult_52_n650), .ZN(mult_52_n417) );
  XNOR2_X1 mult_52_U428 ( .A(B2[3]), .B(n158), .ZN(mult_52_n649) );
  OAI22_X1 mult_52_U427 ( .A1(mult_52_n649), .A2(mult_52_n648), .B1(
        mult_52_n651), .B2(mult_52_n650), .ZN(mult_52_n418) );
  OAI22_X1 mult_52_U426 ( .A1(mult_52_n647), .A2(mult_52_n648), .B1(
        mult_52_n649), .B2(mult_52_n650), .ZN(mult_52_n419) );
  OAI21_X1 mult_52_U425 ( .B1(mult_52_n644), .B2(mult_52_n645), .A(
        mult_52_n646), .ZN(mult_52_n643) );
  XOR2_X1 mult_52_U424 ( .A(mult_52_n643), .B(mult_52_n136), .Z(mult_52_n642)
         );
  XNOR2_X1 mult_52_U423 ( .A(mult_52_n162), .B(mult_52_n642), .ZN(temp4_26_)
         );
  INV_X1 mult_52_U422 ( .A(n168), .ZN(mult_52_n640) );
  INV_X1 mult_52_U421 ( .A(n166), .ZN(mult_52_n639) );
  INV_X1 mult_52_U420 ( .A(n164), .ZN(mult_52_n638) );
  INV_X1 mult_52_U419 ( .A(n162), .ZN(mult_52_n637) );
  XOR2_X2 mult_52_U418 ( .A(reg2[12]), .B(mult_52_n640), .Z(mult_52_n748) );
  XOR2_X2 mult_52_U417 ( .A(reg2[10]), .B(mult_52_n639), .Z(mult_52_n731) );
  XOR2_X2 mult_52_U416 ( .A(reg2[8]), .B(mult_52_n638), .Z(mult_52_n714) );
  XOR2_X2 mult_52_U415 ( .A(reg2[6]), .B(mult_52_n637), .Z(mult_52_n697) );
  XOR2_X2 mult_52_U414 ( .A(reg2[4]), .B(mult_52_n636), .Z(mult_52_n680) );
  INV_X1 mult_52_U413 ( .A(reg2[0]), .ZN(mult_52_n650) );
  INV_X1 mult_52_U412 ( .A(mult_52_n798), .ZN(mult_52_n664) );
  INV_X1 mult_52_U411 ( .A(n170), .ZN(mult_52_n641) );
  INV_X1 mult_52_U410 ( .A(n160), .ZN(mult_52_n636) );
  INV_X1 mult_52_U409 ( .A(n158), .ZN(mult_52_n635) );
  HA_X1 mult_52_U145 ( .A(mult_52_n406), .B(mult_52_n419), .CO(mult_52_n315), 
        .S(mult_52_n316) );
  FA_X1 mult_52_U144 ( .A(mult_52_n418), .B(mult_52_n393), .CI(mult_52_n405), 
        .CO(mult_52_n313), .S(mult_52_n314) );
  HA_X1 mult_52_U143 ( .A(mult_52_n321), .B(mult_52_n392), .CO(mult_52_n311), 
        .S(mult_52_n312) );
  FA_X1 mult_52_U142 ( .A(mult_52_n404), .B(mult_52_n417), .CI(mult_52_n312), 
        .CO(mult_52_n309), .S(mult_52_n310) );
  FA_X1 mult_52_U141 ( .A(mult_52_n416), .B(mult_52_n379), .CI(mult_52_n403), 
        .CO(mult_52_n307), .S(mult_52_n308) );
  FA_X1 mult_52_U140 ( .A(mult_52_n311), .B(mult_52_n391), .CI(mult_52_n308), 
        .CO(mult_52_n305), .S(mult_52_n306) );
  HA_X1 mult_52_U139 ( .A(mult_52_n320), .B(mult_52_n378), .CO(mult_52_n303), 
        .S(mult_52_n304) );
  FA_X1 mult_52_U138 ( .A(mult_52_n390), .B(mult_52_n415), .CI(mult_52_n402), 
        .CO(mult_52_n301), .S(mult_52_n302) );
  FA_X1 mult_52_U137 ( .A(mult_52_n307), .B(mult_52_n304), .CI(mult_52_n302), 
        .CO(mult_52_n299), .S(mult_52_n300) );
  FA_X1 mult_52_U136 ( .A(mult_52_n389), .B(mult_52_n365), .CI(mult_52_n414), 
        .CO(mult_52_n297), .S(mult_52_n298) );
  FA_X1 mult_52_U135 ( .A(mult_52_n377), .B(mult_52_n401), .CI(mult_52_n303), 
        .CO(mult_52_n295), .S(mult_52_n296) );
  FA_X1 mult_52_U134 ( .A(mult_52_n298), .B(mult_52_n301), .CI(mult_52_n296), 
        .CO(mult_52_n293), .S(mult_52_n294) );
  HA_X1 mult_52_U133 ( .A(mult_52_n319), .B(mult_52_n364), .CO(mult_52_n291), 
        .S(mult_52_n292) );
  FA_X1 mult_52_U132 ( .A(mult_52_n376), .B(mult_52_n388), .CI(mult_52_n400), 
        .CO(mult_52_n289), .S(mult_52_n290) );
  FA_X1 mult_52_U131 ( .A(mult_52_n292), .B(mult_52_n413), .CI(mult_52_n297), 
        .CO(mult_52_n287), .S(mult_52_n288) );
  FA_X1 mult_52_U130 ( .A(mult_52_n290), .B(mult_52_n295), .CI(mult_52_n288), 
        .CO(mult_52_n285), .S(mult_52_n286) );
  FA_X1 mult_52_U129 ( .A(mult_52_n375), .B(mult_52_n351), .CI(mult_52_n412), 
        .CO(mult_52_n283), .S(mult_52_n284) );
  FA_X1 mult_52_U128 ( .A(mult_52_n363), .B(mult_52_n399), .CI(mult_52_n387), 
        .CO(mult_52_n281), .S(mult_52_n282) );
  FA_X1 mult_52_U127 ( .A(mult_52_n289), .B(mult_52_n291), .CI(mult_52_n284), 
        .CO(mult_52_n279), .S(mult_52_n280) );
  FA_X1 mult_52_U126 ( .A(mult_52_n287), .B(mult_52_n282), .CI(mult_52_n280), 
        .CO(mult_52_n277), .S(mult_52_n278) );
  HA_X1 mult_52_U125 ( .A(mult_52_n318), .B(mult_52_n350), .CO(mult_52_n275), 
        .S(mult_52_n276) );
  FA_X1 mult_52_U124 ( .A(mult_52_n362), .B(mult_52_n386), .CI(mult_52_n411), 
        .CO(mult_52_n273), .S(mult_52_n274) );
  FA_X1 mult_52_U123 ( .A(mult_52_n374), .B(mult_52_n398), .CI(mult_52_n276), 
        .CO(mult_52_n271), .S(mult_52_n272) );
  FA_X1 mult_52_U122 ( .A(mult_52_n281), .B(mult_52_n283), .CI(mult_52_n274), 
        .CO(mult_52_n269), .S(mult_52_n270) );
  FA_X1 mult_52_U121 ( .A(mult_52_n279), .B(mult_52_n272), .CI(mult_52_n270), 
        .CO(mult_52_n267), .S(mult_52_n268) );
  FA_X1 mult_52_U120 ( .A(mult_52_n361), .B(mult_52_n337), .CI(mult_52_n410), 
        .CO(mult_52_n265), .S(mult_52_n266) );
  FA_X1 mult_52_U109 ( .A(mult_52_n349), .B(mult_52_n397), .CI(mult_52_n373), 
        .CO(mult_52_n263), .S(mult_52_n264) );
  FA_X1 mult_52_U108 ( .A(mult_52_n275), .B(mult_52_n385), .CI(mult_52_n273), 
        .CO(mult_52_n261), .S(mult_52_n262) );
  FA_X1 mult_52_U107 ( .A(mult_52_n264), .B(mult_52_n266), .CI(mult_52_n271), 
        .CO(mult_52_n259), .S(mult_52_n260) );
  FA_X1 mult_52_U106 ( .A(mult_52_n262), .B(mult_52_n269), .CI(mult_52_n260), 
        .CO(mult_52_n257), .S(mult_52_n258) );
  HA_X1 mult_52_U105 ( .A(mult_52_n317), .B(mult_52_n336), .CO(mult_52_n255), 
        .S(mult_52_n256) );
  FA_X1 mult_52_U104 ( .A(mult_52_n409), .B(mult_52_n372), .CI(mult_52_n396), 
        .CO(mult_52_n253), .S(mult_52_n254) );
  FA_X1 mult_52_U103 ( .A(mult_52_n348), .B(mult_52_n384), .CI(mult_52_n360), 
        .CO(mult_52_n251), .S(mult_52_n252) );
  FA_X1 mult_52_U102 ( .A(mult_52_n265), .B(mult_52_n256), .CI(mult_52_n263), 
        .CO(mult_52_n249), .S(mult_52_n250) );
  FA_X1 mult_52_U101 ( .A(mult_52_n254), .B(mult_52_n252), .CI(mult_52_n261), 
        .CO(mult_52_n247), .S(mult_52_n248) );
  FA_X1 mult_52_U100 ( .A(mult_52_n259), .B(mult_52_n250), .CI(mult_52_n248), 
        .CO(mult_52_n245), .S(mult_52_n246) );
  FA_X1 mult_52_U97 ( .A(mult_52_n395), .B(mult_52_n359), .CI(mult_52_n408), 
        .CO(mult_52_n241), .S(mult_52_n242) );
  FA_X1 mult_52_U96 ( .A(mult_52_n335), .B(mult_52_n371), .CI(mult_52_n255), 
        .CO(mult_52_n239), .S(mult_52_n240) );
  FA_X1 mult_52_U95 ( .A(mult_52_n253), .B(mult_52_n244), .CI(mult_52_n251), 
        .CO(mult_52_n237), .S(mult_52_n238) );
  FA_X1 mult_52_U94 ( .A(mult_52_n240), .B(mult_52_n242), .CI(mult_52_n249), 
        .CO(mult_52_n235), .S(mult_52_n236) );
  FA_X1 mult_52_U93 ( .A(mult_52_n247), .B(mult_52_n238), .CI(mult_52_n236), 
        .CO(mult_52_n233), .S(mult_52_n234) );
  FA_X1 mult_52_U91 ( .A(mult_52_n382), .B(mult_52_n346), .CI(mult_52_n232), 
        .CO(mult_52_n229), .S(mult_52_n230) );
  FA_X1 mult_52_U90 ( .A(mult_52_n334), .B(mult_52_n370), .CI(mult_52_n358), 
        .CO(mult_52_n227), .S(mult_52_n228) );
  FA_X1 mult_52_U89 ( .A(mult_52_n241), .B(mult_52_n243), .CI(mult_52_n239), 
        .CO(mult_52_n225), .S(mult_52_n226) );
  FA_X1 mult_52_U88 ( .A(mult_52_n230), .B(mult_52_n228), .CI(mult_52_n237), 
        .CO(mult_52_n223), .S(mult_52_n224) );
  FA_X1 mult_52_U87 ( .A(mult_52_n235), .B(mult_52_n226), .CI(mult_52_n224), 
        .CO(mult_52_n221), .S(mult_52_n222) );
  FA_X1 mult_52_U86 ( .A(mult_52_n231), .B(mult_52_n333), .CI(mult_52_n394), 
        .CO(mult_52_n219), .S(mult_52_n220) );
  FA_X1 mult_52_U85 ( .A(mult_52_n345), .B(mult_52_n381), .CI(mult_52_n357), 
        .CO(mult_52_n217), .S(mult_52_n218) );
  FA_X1 mult_52_U84 ( .A(mult_52_n229), .B(mult_52_n369), .CI(mult_52_n227), 
        .CO(mult_52_n215), .S(mult_52_n216) );
  FA_X1 mult_52_U83 ( .A(mult_52_n220), .B(mult_52_n218), .CI(mult_52_n225), 
        .CO(mult_52_n213), .S(mult_52_n214) );
  FA_X1 mult_52_U82 ( .A(mult_52_n223), .B(mult_52_n216), .CI(mult_52_n214), 
        .CO(mult_52_n211), .S(mult_52_n212) );
  FA_X1 mult_52_U80 ( .A(mult_52_n368), .B(mult_52_n344), .CI(mult_52_n210), 
        .CO(mult_52_n207), .S(mult_52_n208) );
  FA_X1 mult_52_U79 ( .A(mult_52_n332), .B(mult_52_n356), .CI(mult_52_n219), 
        .CO(mult_52_n205), .S(mult_52_n206) );
  FA_X1 mult_52_U78 ( .A(mult_52_n208), .B(mult_52_n217), .CI(mult_52_n215), 
        .CO(mult_52_n203), .S(mult_52_n204) );
  FA_X1 mult_52_U77 ( .A(mult_52_n213), .B(mult_52_n206), .CI(mult_52_n204), 
        .CO(mult_52_n201), .S(mult_52_n202) );
  FA_X1 mult_52_U76 ( .A(mult_52_n209), .B(mult_52_n331), .CI(mult_52_n380), 
        .CO(mult_52_n199), .S(mult_52_n200) );
  FA_X1 mult_52_U75 ( .A(mult_52_n355), .B(mult_52_n343), .CI(mult_52_n367), 
        .CO(mult_52_n197), .S(mult_52_n198) );
  FA_X1 mult_52_U74 ( .A(mult_52_n198), .B(mult_52_n207), .CI(mult_52_n200), 
        .CO(mult_52_n195), .S(mult_52_n196) );
  FA_X1 mult_52_U73 ( .A(mult_52_n203), .B(mult_52_n205), .CI(mult_52_n196), 
        .CO(mult_52_n193), .S(mult_52_n194) );
  FA_X1 mult_52_U71 ( .A(mult_52_n330), .B(mult_52_n342), .CI(mult_52_n192), 
        .CO(mult_52_n189), .S(mult_52_n190) );
  FA_X1 mult_52_U70 ( .A(mult_52_n199), .B(mult_52_n354), .CI(mult_52_n197), 
        .CO(mult_52_n187), .S(mult_52_n188) );
  FA_X1 mult_52_U69 ( .A(mult_52_n188), .B(mult_52_n190), .CI(mult_52_n195), 
        .CO(mult_52_n185), .S(mult_52_n186) );
  FA_X1 mult_52_U68 ( .A(mult_52_n191), .B(mult_52_n329), .CI(mult_52_n366), 
        .CO(mult_52_n183), .S(mult_52_n184) );
  FA_X1 mult_52_U67 ( .A(mult_52_n341), .B(mult_52_n353), .CI(mult_52_n189), 
        .CO(mult_52_n181), .S(mult_52_n182) );
  FA_X1 mult_52_U66 ( .A(mult_52_n187), .B(mult_52_n184), .CI(mult_52_n182), 
        .CO(mult_52_n179), .S(mult_52_n180) );
  FA_X1 mult_52_U64 ( .A(mult_52_n328), .B(mult_52_n340), .CI(mult_52_n178), 
        .CO(mult_52_n175), .S(mult_52_n176) );
  FA_X1 mult_52_U63 ( .A(mult_52_n176), .B(mult_52_n183), .CI(mult_52_n181), 
        .CO(mult_52_n173), .S(mult_52_n174) );
  FA_X1 mult_52_U62 ( .A(mult_52_n327), .B(mult_52_n177), .CI(mult_52_n352), 
        .CO(mult_52_n171), .S(mult_52_n172) );
  FA_X1 mult_52_U61 ( .A(mult_52_n175), .B(mult_52_n339), .CI(mult_52_n172), 
        .CO(mult_52_n169), .S(mult_52_n170) );
  FA_X1 mult_52_U59 ( .A(mult_52_n168), .B(mult_52_n326), .CI(mult_52_n171), 
        .CO(mult_52_n165), .S(mult_52_n166) );
  FA_X1 mult_52_U58 ( .A(mult_52_n325), .B(mult_52_n167), .CI(mult_52_n338), 
        .CO(mult_52_n163), .S(mult_52_n164) );
  FA_X1 mult_52_U44 ( .A(mult_52_n246), .B(mult_52_n257), .CI(mult_52_n149), 
        .CO(mult_52_n148), .S(temp4_13_) );
  FA_X1 mult_52_U43 ( .A(mult_52_n234), .B(mult_52_n245), .CI(mult_52_n148), 
        .CO(mult_52_n147), .S(temp4_14_) );
  FA_X1 mult_52_U42 ( .A(mult_52_n222), .B(mult_52_n233), .CI(mult_52_n147), 
        .CO(mult_52_n146), .S(temp4_15_) );
  FA_X1 mult_52_U41 ( .A(mult_52_n212), .B(mult_52_n221), .CI(mult_52_n146), 
        .CO(mult_52_n145), .S(temp4_16_) );
  FA_X1 mult_52_U40 ( .A(mult_52_n202), .B(mult_52_n211), .CI(mult_52_n145), 
        .CO(mult_52_n144), .S(temp4_17_) );
  FA_X1 mult_52_U39 ( .A(mult_52_n194), .B(mult_52_n201), .CI(mult_52_n144), 
        .CO(mult_52_n143), .S(temp4_18_) );
  FA_X1 mult_52_U38 ( .A(mult_52_n186), .B(mult_52_n193), .CI(mult_52_n143), 
        .CO(mult_52_n142), .S(temp4_19_) );
  FA_X1 mult_52_U37 ( .A(mult_52_n180), .B(mult_52_n185), .CI(mult_52_n142), 
        .CO(mult_52_n141), .S(temp4_20_) );
  FA_X1 mult_52_U30 ( .A(mult_52_n174), .B(mult_52_n179), .CI(mult_52_n141), 
        .CO(mult_52_n140), .S(temp4_21_) );
  FA_X1 mult_52_U20 ( .A(mult_52_n170), .B(mult_52_n173), .CI(mult_52_n140), 
        .CO(mult_52_n139), .S(temp4_22_) );
  FA_X1 mult_52_U10 ( .A(mult_52_n166), .B(mult_52_n169), .CI(mult_52_n139), 
        .CO(mult_52_n138), .S(temp4_23_) );
  FA_X1 mult_52_U9 ( .A(mult_52_n165), .B(mult_52_n164), .CI(mult_52_n138), 
        .CO(mult_52_n137), .S(temp4_24_) );
  FA_X1 mult_52_U8 ( .A(mult_52_n163), .B(mult_52_n162), .CI(mult_52_n137), 
        .CO(mult_52_n136), .S(temp4_25_) );
  XOR2_X1 add_1_root_add_0_root_add_59_U2 ( .A(temp3_13_), .B(temp4_13_), .Z(
        ff_0_) );
  AND2_X1 add_1_root_add_0_root_add_59_U1 ( .A1(temp4_13_), .A2(temp3_13_), 
        .ZN(add_1_root_add_0_root_add_59_carry_1_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_1 ( .A(temp4_14_), .B(temp3_14_), .CI(
        add_1_root_add_0_root_add_59_carry_1_), .CO(
        add_1_root_add_0_root_add_59_carry_2_), .S(ff_1_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_2 ( .A(temp4_15_), .B(temp3_15_), .CI(
        add_1_root_add_0_root_add_59_carry_2_), .CO(
        add_1_root_add_0_root_add_59_carry_3_), .S(ff_2_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_3 ( .A(temp4_16_), .B(temp3_16_), .CI(
        add_1_root_add_0_root_add_59_carry_3_), .CO(
        add_1_root_add_0_root_add_59_carry_4_), .S(ff_3_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_4 ( .A(temp4_17_), .B(temp3_17_), .CI(
        add_1_root_add_0_root_add_59_carry_4_), .CO(
        add_1_root_add_0_root_add_59_carry_5_), .S(ff_4_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_5 ( .A(temp4_18_), .B(temp3_18_), .CI(
        add_1_root_add_0_root_add_59_carry_5_), .CO(
        add_1_root_add_0_root_add_59_carry_6_), .S(ff_5_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_6 ( .A(temp4_19_), .B(temp3_19_), .CI(
        add_1_root_add_0_root_add_59_carry_6_), .CO(
        add_1_root_add_0_root_add_59_carry_7_), .S(ff_6_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_7 ( .A(temp4_20_), .B(temp3_20_), .CI(
        add_1_root_add_0_root_add_59_carry_7_), .CO(
        add_1_root_add_0_root_add_59_carry_8_), .S(ff_7_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_8 ( .A(temp4_21_), .B(temp3_21_), .CI(
        add_1_root_add_0_root_add_59_carry_8_), .CO(
        add_1_root_add_0_root_add_59_carry_9_), .S(ff_8_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_9 ( .A(temp4_22_), .B(temp3_22_), .CI(
        add_1_root_add_0_root_add_59_carry_9_), .CO(
        add_1_root_add_0_root_add_59_carry_10_), .S(ff_9_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_10 ( .A(temp4_23_), .B(temp3_23_), 
        .CI(add_1_root_add_0_root_add_59_carry_10_), .CO(
        add_1_root_add_0_root_add_59_carry_11_), .S(ff_10_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_11 ( .A(temp4_24_), .B(temp3_24_), 
        .CI(add_1_root_add_0_root_add_59_carry_11_), .CO(
        add_1_root_add_0_root_add_59_carry_12_), .S(ff_11_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_12 ( .A(temp4_25_), .B(temp3_25_), 
        .CI(add_1_root_add_0_root_add_59_carry_12_), .CO(
        add_1_root_add_0_root_add_59_carry_13_), .S(ff_12_) );
  FA_X1 add_1_root_add_0_root_add_59_U1_13 ( .A(temp4_26_), .B(temp3_26_), 
        .CI(add_1_root_add_0_root_add_59_carry_13_), .S(ff_13_) );
  XOR2_X1 mult_54_U691 ( .A(w[2]), .B(w[1]), .Z(mult_54_n798) );
  INV_X1 mult_54_U690 ( .A(w[1]), .ZN(mult_54_n655) );
  NOR2_X1 mult_54_U689 ( .A1(mult_54_n655), .A2(B0[1]), .ZN(mult_54_n803) );
  INV_X1 mult_54_U688 ( .A(mult_54_n803), .ZN(mult_54_n805) );
  NAND2_X1 mult_54_U687 ( .A1(w[1]), .A2(mult_54_n643), .ZN(mult_54_n641) );
  XNOR2_X1 mult_54_U686 ( .A(B0[2]), .B(w[1]), .ZN(mult_54_n640) );
  OAI22_X1 mult_54_U685 ( .A1(mult_54_n805), .A2(mult_54_n641), .B1(
        mult_54_n640), .B2(mult_54_n643), .ZN(mult_54_n804) );
  NAND2_X1 mult_54_U684 ( .A1(mult_54_n798), .A2(mult_54_n804), .ZN(
        mult_54_n801) );
  NAND2_X1 mult_54_U683 ( .A1(mult_54_n803), .A2(mult_54_n804), .ZN(
        mult_54_n802) );
  INV_X1 mult_54_U682 ( .A(B0[0]), .ZN(mult_54_n673) );
  MUX2_X1 mult_54_U681 ( .A(mult_54_n801), .B(mult_54_n802), .S(mult_54_n673), 
        .Z(mult_54_n800) );
  INV_X1 mult_54_U680 ( .A(mult_54_n800), .ZN(mult_54_n795) );
  INV_X1 mult_54_U679 ( .A(w[3]), .ZN(mult_54_n771) );
  XNOR2_X1 mult_54_U678 ( .A(mult_54_n771), .B(w[2]), .ZN(mult_54_n799) );
  NAND2_X1 mult_54_U677 ( .A1(mult_54_n658), .A2(mult_54_n799), .ZN(
        mult_54_n657) );
  NAND3_X1 mult_54_U676 ( .A1(mult_54_n798), .A2(mult_54_n673), .A3(w[3]), 
        .ZN(mult_54_n797) );
  OAI21_X1 mult_54_U675 ( .B1(mult_54_n771), .B2(mult_54_n657), .A(
        mult_54_n797), .ZN(mult_54_n796) );
  AOI222_X1 mult_54_U674 ( .A1(mult_54_n795), .A2(mult_54_n316), .B1(
        mult_54_n796), .B2(mult_54_n795), .C1(mult_54_n796), .C2(mult_54_n316), 
        .ZN(mult_54_n794) );
  INV_X1 mult_54_U673 ( .A(mult_54_n794), .ZN(mult_54_n793) );
  AOI222_X1 mult_54_U672 ( .A1(mult_54_n793), .A2(mult_54_n314), .B1(
        mult_54_n793), .B2(mult_54_n315), .C1(mult_54_n315), .C2(mult_54_n314), 
        .ZN(mult_54_n792) );
  INV_X1 mult_54_U671 ( .A(mult_54_n792), .ZN(mult_54_n791) );
  AOI222_X1 mult_54_U670 ( .A1(mult_54_n791), .A2(mult_54_n310), .B1(
        mult_54_n791), .B2(mult_54_n313), .C1(mult_54_n313), .C2(mult_54_n310), 
        .ZN(mult_54_n790) );
  INV_X1 mult_54_U669 ( .A(mult_54_n790), .ZN(mult_54_n789) );
  AOI222_X1 mult_54_U668 ( .A1(mult_54_n789), .A2(mult_54_n306), .B1(
        mult_54_n789), .B2(mult_54_n309), .C1(mult_54_n309), .C2(mult_54_n306), 
        .ZN(mult_54_n788) );
  INV_X1 mult_54_U667 ( .A(mult_54_n788), .ZN(mult_54_n787) );
  AOI222_X1 mult_54_U666 ( .A1(mult_54_n787), .A2(mult_54_n300), .B1(
        mult_54_n787), .B2(mult_54_n305), .C1(mult_54_n305), .C2(mult_54_n300), 
        .ZN(mult_54_n786) );
  INV_X1 mult_54_U665 ( .A(mult_54_n786), .ZN(mult_54_n785) );
  AOI222_X1 mult_54_U664 ( .A1(mult_54_n785), .A2(mult_54_n294), .B1(
        mult_54_n785), .B2(mult_54_n299), .C1(mult_54_n299), .C2(mult_54_n294), 
        .ZN(mult_54_n784) );
  INV_X1 mult_54_U663 ( .A(mult_54_n784), .ZN(mult_54_n783) );
  AOI222_X1 mult_54_U662 ( .A1(mult_54_n783), .A2(mult_54_n286), .B1(
        mult_54_n783), .B2(mult_54_n293), .C1(mult_54_n293), .C2(mult_54_n286), 
        .ZN(mult_54_n780) );
  INV_X1 mult_54_U661 ( .A(mult_54_n278), .ZN(mult_54_n781) );
  INV_X1 mult_54_U660 ( .A(mult_54_n285), .ZN(mult_54_n782) );
  OAI222_X1 mult_54_U659 ( .A1(mult_54_n780), .A2(mult_54_n781), .B1(
        mult_54_n780), .B2(mult_54_n782), .C1(mult_54_n782), .C2(mult_54_n781), 
        .ZN(mult_54_n779) );
  AOI222_X1 mult_54_U658 ( .A1(mult_54_n779), .A2(mult_54_n268), .B1(
        mult_54_n779), .B2(mult_54_n277), .C1(mult_54_n277), .C2(mult_54_n268), 
        .ZN(mult_54_n776) );
  INV_X1 mult_54_U657 ( .A(mult_54_n258), .ZN(mult_54_n777) );
  INV_X1 mult_54_U656 ( .A(mult_54_n267), .ZN(mult_54_n778) );
  OAI222_X1 mult_54_U655 ( .A1(mult_54_n776), .A2(mult_54_n777), .B1(
        mult_54_n776), .B2(mult_54_n778), .C1(mult_54_n778), .C2(mult_54_n777), 
        .ZN(mult_54_n149) );
  XOR2_X1 mult_54_U654 ( .A(B0[12]), .B(w[13]), .Z(mult_54_n757) );
  INV_X1 mult_54_U653 ( .A(w[11]), .ZN(mult_54_n764) );
  INV_X1 mult_54_U652 ( .A(w[13]), .ZN(mult_54_n766) );
  XNOR2_X1 mult_54_U651 ( .A(mult_54_n766), .B(w[12]), .ZN(mult_54_n775) );
  NAND2_X1 mult_54_U650 ( .A1(mult_54_n742), .A2(mult_54_n775), .ZN(
        mult_54_n744) );
  INV_X1 mult_54_U649 ( .A(mult_54_n744), .ZN(mult_54_n637) );
  INV_X1 mult_54_U648 ( .A(mult_54_n742), .ZN(mult_54_n638) );
  XNOR2_X1 mult_54_U647 ( .A(B0[13]), .B(mult_54_n766), .ZN(mult_54_n639) );
  AOI22_X1 mult_54_U646 ( .A1(mult_54_n757), .A2(mult_54_n637), .B1(
        mult_54_n638), .B2(mult_54_n639), .ZN(mult_54_n162) );
  XNOR2_X1 mult_54_U645 ( .A(B0[12]), .B(w[11]), .ZN(mult_54_n739) );
  INV_X1 mult_54_U644 ( .A(w[9]), .ZN(mult_54_n762) );
  XNOR2_X1 mult_54_U643 ( .A(mult_54_n764), .B(w[10]), .ZN(mult_54_n774) );
  NAND2_X1 mult_54_U642 ( .A1(mult_54_n725), .A2(mult_54_n774), .ZN(
        mult_54_n727) );
  XNOR2_X1 mult_54_U641 ( .A(B0[13]), .B(w[11]), .ZN(mult_54_n741) );
  OAI22_X1 mult_54_U640 ( .A1(mult_54_n739), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n741), .ZN(mult_54_n167) );
  INV_X1 mult_54_U639 ( .A(mult_54_n167), .ZN(mult_54_n168) );
  XNOR2_X1 mult_54_U638 ( .A(B0[12]), .B(w[9]), .ZN(mult_54_n722) );
  INV_X1 mult_54_U637 ( .A(w[7]), .ZN(mult_54_n760) );
  XNOR2_X1 mult_54_U636 ( .A(mult_54_n762), .B(w[8]), .ZN(mult_54_n773) );
  NAND2_X1 mult_54_U635 ( .A1(mult_54_n708), .A2(mult_54_n773), .ZN(
        mult_54_n710) );
  XNOR2_X1 mult_54_U634 ( .A(B0[13]), .B(w[9]), .ZN(mult_54_n724) );
  OAI22_X1 mult_54_U633 ( .A1(mult_54_n722), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n724), .ZN(mult_54_n177) );
  INV_X1 mult_54_U632 ( .A(mult_54_n177), .ZN(mult_54_n178) );
  XNOR2_X1 mult_54_U631 ( .A(B0[12]), .B(w[7]), .ZN(mult_54_n705) );
  INV_X1 mult_54_U630 ( .A(w[5]), .ZN(mult_54_n758) );
  XNOR2_X1 mult_54_U629 ( .A(mult_54_n760), .B(w[6]), .ZN(mult_54_n772) );
  NAND2_X1 mult_54_U628 ( .A1(mult_54_n691), .A2(mult_54_n772), .ZN(
        mult_54_n693) );
  XNOR2_X1 mult_54_U627 ( .A(B0[13]), .B(w[7]), .ZN(mult_54_n707) );
  OAI22_X1 mult_54_U626 ( .A1(mult_54_n705), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n707), .ZN(mult_54_n191) );
  INV_X1 mult_54_U625 ( .A(mult_54_n191), .ZN(mult_54_n192) );
  XNOR2_X1 mult_54_U624 ( .A(B0[12]), .B(w[5]), .ZN(mult_54_n688) );
  XNOR2_X1 mult_54_U623 ( .A(mult_54_n758), .B(w[4]), .ZN(mult_54_n770) );
  NAND2_X1 mult_54_U622 ( .A1(mult_54_n674), .A2(mult_54_n770), .ZN(
        mult_54_n676) );
  XNOR2_X1 mult_54_U621 ( .A(B0[13]), .B(w[5]), .ZN(mult_54_n690) );
  OAI22_X1 mult_54_U620 ( .A1(mult_54_n688), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n690), .ZN(mult_54_n209) );
  INV_X1 mult_54_U619 ( .A(mult_54_n209), .ZN(mult_54_n210) );
  XNOR2_X1 mult_54_U618 ( .A(B0[12]), .B(w[3]), .ZN(mult_54_n670) );
  XNOR2_X1 mult_54_U617 ( .A(B0[13]), .B(w[3]), .ZN(mult_54_n672) );
  OAI22_X1 mult_54_U616 ( .A1(mult_54_n670), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n672), .ZN(mult_54_n231) );
  INV_X1 mult_54_U615 ( .A(mult_54_n231), .ZN(mult_54_n232) );
  XNOR2_X1 mult_54_U614 ( .A(B0[3]), .B(w[11]), .ZN(mult_54_n730) );
  XNOR2_X1 mult_54_U613 ( .A(B0[4]), .B(w[11]), .ZN(mult_54_n731) );
  OAI22_X1 mult_54_U612 ( .A1(mult_54_n730), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n731), .ZN(mult_54_n768) );
  XNOR2_X1 mult_54_U611 ( .A(B0[9]), .B(w[5]), .ZN(mult_54_n685) );
  XNOR2_X1 mult_54_U610 ( .A(B0[10]), .B(w[5]), .ZN(mult_54_n686) );
  OAI22_X1 mult_54_U609 ( .A1(mult_54_n685), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n686), .ZN(mult_54_n769) );
  OR2_X1 mult_54_U608 ( .A1(mult_54_n768), .A2(mult_54_n769), .ZN(mult_54_n243) );
  XNOR2_X1 mult_54_U607 ( .A(mult_54_n768), .B(mult_54_n769), .ZN(mult_54_n244) );
  NAND3_X1 mult_54_U606 ( .A1(mult_54_n638), .A2(mult_54_n673), .A3(w[13]), 
        .ZN(mult_54_n767) );
  OAI21_X1 mult_54_U605 ( .B1(mult_54_n766), .B2(mult_54_n744), .A(
        mult_54_n767), .ZN(mult_54_n317) );
  OR3_X1 mult_54_U604 ( .A1(mult_54_n725), .A2(B0[0]), .A3(mult_54_n764), .ZN(
        mult_54_n765) );
  OAI21_X1 mult_54_U603 ( .B1(mult_54_n764), .B2(mult_54_n727), .A(
        mult_54_n765), .ZN(mult_54_n318) );
  OR3_X1 mult_54_U602 ( .A1(mult_54_n708), .A2(B0[0]), .A3(mult_54_n762), .ZN(
        mult_54_n763) );
  OAI21_X1 mult_54_U601 ( .B1(mult_54_n762), .B2(mult_54_n710), .A(
        mult_54_n763), .ZN(mult_54_n319) );
  OR3_X1 mult_54_U600 ( .A1(mult_54_n691), .A2(B0[0]), .A3(mult_54_n760), .ZN(
        mult_54_n761) );
  OAI21_X1 mult_54_U599 ( .B1(mult_54_n760), .B2(mult_54_n693), .A(
        mult_54_n761), .ZN(mult_54_n320) );
  OR3_X1 mult_54_U598 ( .A1(mult_54_n674), .A2(B0[0]), .A3(mult_54_n758), .ZN(
        mult_54_n759) );
  OAI21_X1 mult_54_U597 ( .B1(mult_54_n758), .B2(mult_54_n676), .A(
        mult_54_n759), .ZN(mult_54_n321) );
  XNOR2_X1 mult_54_U596 ( .A(B0[11]), .B(w[13]), .ZN(mult_54_n755) );
  INV_X1 mult_54_U595 ( .A(mult_54_n757), .ZN(mult_54_n756) );
  OAI22_X1 mult_54_U594 ( .A1(mult_54_n755), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n756), .ZN(mult_54_n325) );
  XNOR2_X1 mult_54_U593 ( .A(B0[10]), .B(w[13]), .ZN(mult_54_n754) );
  OAI22_X1 mult_54_U592 ( .A1(mult_54_n754), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n755), .ZN(mult_54_n326) );
  XNOR2_X1 mult_54_U591 ( .A(B0[9]), .B(w[13]), .ZN(mult_54_n753) );
  OAI22_X1 mult_54_U590 ( .A1(mult_54_n753), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n754), .ZN(mult_54_n327) );
  XNOR2_X1 mult_54_U589 ( .A(B0[8]), .B(w[13]), .ZN(mult_54_n752) );
  OAI22_X1 mult_54_U588 ( .A1(mult_54_n752), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n753), .ZN(mult_54_n328) );
  XNOR2_X1 mult_54_U587 ( .A(B0[7]), .B(w[13]), .ZN(mult_54_n751) );
  OAI22_X1 mult_54_U586 ( .A1(mult_54_n751), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n752), .ZN(mult_54_n329) );
  XNOR2_X1 mult_54_U585 ( .A(B0[6]), .B(w[13]), .ZN(mult_54_n750) );
  OAI22_X1 mult_54_U584 ( .A1(mult_54_n750), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n751), .ZN(mult_54_n330) );
  XNOR2_X1 mult_54_U583 ( .A(B0[5]), .B(w[13]), .ZN(mult_54_n749) );
  OAI22_X1 mult_54_U582 ( .A1(mult_54_n749), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n750), .ZN(mult_54_n331) );
  XNOR2_X1 mult_54_U581 ( .A(B0[4]), .B(w[13]), .ZN(mult_54_n748) );
  OAI22_X1 mult_54_U580 ( .A1(mult_54_n748), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n749), .ZN(mult_54_n332) );
  XNOR2_X1 mult_54_U579 ( .A(B0[3]), .B(w[13]), .ZN(mult_54_n747) );
  OAI22_X1 mult_54_U578 ( .A1(mult_54_n747), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n748), .ZN(mult_54_n333) );
  XNOR2_X1 mult_54_U577 ( .A(B0[2]), .B(w[13]), .ZN(mult_54_n746) );
  OAI22_X1 mult_54_U576 ( .A1(mult_54_n746), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n747), .ZN(mult_54_n334) );
  XNOR2_X1 mult_54_U575 ( .A(B0[1]), .B(w[13]), .ZN(mult_54_n745) );
  OAI22_X1 mult_54_U574 ( .A1(mult_54_n745), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n746), .ZN(mult_54_n335) );
  XNOR2_X1 mult_54_U573 ( .A(w[13]), .B(B0[0]), .ZN(mult_54_n743) );
  OAI22_X1 mult_54_U572 ( .A1(mult_54_n743), .A2(mult_54_n744), .B1(
        mult_54_n742), .B2(mult_54_n745), .ZN(mult_54_n336) );
  NOR2_X1 mult_54_U571 ( .A1(mult_54_n673), .A2(mult_54_n742), .ZN(
        mult_54_n337) );
  AOI21_X1 mult_54_U570 ( .B1(mult_54_n727), .B2(mult_54_n725), .A(
        mult_54_n741), .ZN(mult_54_n740) );
  INV_X1 mult_54_U569 ( .A(mult_54_n740), .ZN(mult_54_n338) );
  XNOR2_X1 mult_54_U568 ( .A(B0[11]), .B(w[11]), .ZN(mult_54_n738) );
  OAI22_X1 mult_54_U567 ( .A1(mult_54_n738), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n739), .ZN(mult_54_n339) );
  XNOR2_X1 mult_54_U566 ( .A(B0[10]), .B(w[11]), .ZN(mult_54_n737) );
  OAI22_X1 mult_54_U565 ( .A1(mult_54_n737), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n738), .ZN(mult_54_n340) );
  XNOR2_X1 mult_54_U564 ( .A(B0[9]), .B(w[11]), .ZN(mult_54_n736) );
  OAI22_X1 mult_54_U563 ( .A1(mult_54_n736), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n737), .ZN(mult_54_n341) );
  XNOR2_X1 mult_54_U562 ( .A(B0[8]), .B(w[11]), .ZN(mult_54_n735) );
  OAI22_X1 mult_54_U561 ( .A1(mult_54_n735), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n736), .ZN(mult_54_n342) );
  XNOR2_X1 mult_54_U560 ( .A(B0[7]), .B(w[11]), .ZN(mult_54_n734) );
  OAI22_X1 mult_54_U559 ( .A1(mult_54_n734), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n735), .ZN(mult_54_n343) );
  XNOR2_X1 mult_54_U558 ( .A(B0[6]), .B(w[11]), .ZN(mult_54_n733) );
  OAI22_X1 mult_54_U557 ( .A1(mult_54_n733), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n734), .ZN(mult_54_n344) );
  XNOR2_X1 mult_54_U556 ( .A(B0[5]), .B(w[11]), .ZN(mult_54_n732) );
  OAI22_X1 mult_54_U555 ( .A1(mult_54_n732), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n733), .ZN(mult_54_n345) );
  OAI22_X1 mult_54_U554 ( .A1(mult_54_n731), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n732), .ZN(mult_54_n346) );
  XNOR2_X1 mult_54_U553 ( .A(B0[2]), .B(w[11]), .ZN(mult_54_n729) );
  OAI22_X1 mult_54_U552 ( .A1(mult_54_n729), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n730), .ZN(mult_54_n348) );
  XNOR2_X1 mult_54_U551 ( .A(B0[1]), .B(w[11]), .ZN(mult_54_n728) );
  OAI22_X1 mult_54_U550 ( .A1(mult_54_n728), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n729), .ZN(mult_54_n349) );
  XNOR2_X1 mult_54_U549 ( .A(w[11]), .B(B0[0]), .ZN(mult_54_n726) );
  OAI22_X1 mult_54_U548 ( .A1(mult_54_n726), .A2(mult_54_n727), .B1(
        mult_54_n725), .B2(mult_54_n728), .ZN(mult_54_n350) );
  NOR2_X1 mult_54_U547 ( .A1(mult_54_n673), .A2(mult_54_n725), .ZN(
        mult_54_n351) );
  AOI21_X1 mult_54_U546 ( .B1(mult_54_n710), .B2(mult_54_n708), .A(
        mult_54_n724), .ZN(mult_54_n723) );
  INV_X1 mult_54_U545 ( .A(mult_54_n723), .ZN(mult_54_n352) );
  XNOR2_X1 mult_54_U544 ( .A(B0[11]), .B(w[9]), .ZN(mult_54_n721) );
  OAI22_X1 mult_54_U543 ( .A1(mult_54_n721), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n722), .ZN(mult_54_n353) );
  XNOR2_X1 mult_54_U542 ( .A(B0[10]), .B(w[9]), .ZN(mult_54_n720) );
  OAI22_X1 mult_54_U541 ( .A1(mult_54_n720), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n721), .ZN(mult_54_n354) );
  XNOR2_X1 mult_54_U540 ( .A(B0[9]), .B(w[9]), .ZN(mult_54_n719) );
  OAI22_X1 mult_54_U539 ( .A1(mult_54_n719), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n720), .ZN(mult_54_n355) );
  XNOR2_X1 mult_54_U538 ( .A(B0[8]), .B(w[9]), .ZN(mult_54_n718) );
  OAI22_X1 mult_54_U537 ( .A1(mult_54_n718), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n719), .ZN(mult_54_n356) );
  XNOR2_X1 mult_54_U536 ( .A(B0[7]), .B(w[9]), .ZN(mult_54_n717) );
  OAI22_X1 mult_54_U535 ( .A1(mult_54_n717), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n718), .ZN(mult_54_n357) );
  XNOR2_X1 mult_54_U534 ( .A(B0[6]), .B(w[9]), .ZN(mult_54_n716) );
  OAI22_X1 mult_54_U533 ( .A1(mult_54_n716), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n717), .ZN(mult_54_n358) );
  XNOR2_X1 mult_54_U532 ( .A(B0[5]), .B(w[9]), .ZN(mult_54_n715) );
  OAI22_X1 mult_54_U531 ( .A1(mult_54_n715), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n716), .ZN(mult_54_n359) );
  XNOR2_X1 mult_54_U530 ( .A(B0[4]), .B(w[9]), .ZN(mult_54_n714) );
  OAI22_X1 mult_54_U529 ( .A1(mult_54_n714), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n715), .ZN(mult_54_n360) );
  XNOR2_X1 mult_54_U528 ( .A(B0[3]), .B(w[9]), .ZN(mult_54_n713) );
  OAI22_X1 mult_54_U527 ( .A1(mult_54_n713), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n714), .ZN(mult_54_n361) );
  XNOR2_X1 mult_54_U526 ( .A(B0[2]), .B(w[9]), .ZN(mult_54_n712) );
  OAI22_X1 mult_54_U525 ( .A1(mult_54_n712), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n713), .ZN(mult_54_n362) );
  XNOR2_X1 mult_54_U524 ( .A(B0[1]), .B(w[9]), .ZN(mult_54_n711) );
  OAI22_X1 mult_54_U523 ( .A1(mult_54_n711), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n712), .ZN(mult_54_n363) );
  XNOR2_X1 mult_54_U522 ( .A(w[9]), .B(B0[0]), .ZN(mult_54_n709) );
  OAI22_X1 mult_54_U521 ( .A1(mult_54_n709), .A2(mult_54_n710), .B1(
        mult_54_n708), .B2(mult_54_n711), .ZN(mult_54_n364) );
  NOR2_X1 mult_54_U520 ( .A1(mult_54_n673), .A2(mult_54_n708), .ZN(
        mult_54_n365) );
  AOI21_X1 mult_54_U519 ( .B1(mult_54_n693), .B2(mult_54_n691), .A(
        mult_54_n707), .ZN(mult_54_n706) );
  INV_X1 mult_54_U518 ( .A(mult_54_n706), .ZN(mult_54_n366) );
  XNOR2_X1 mult_54_U517 ( .A(B0[11]), .B(w[7]), .ZN(mult_54_n704) );
  OAI22_X1 mult_54_U516 ( .A1(mult_54_n704), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n705), .ZN(mult_54_n367) );
  XNOR2_X1 mult_54_U515 ( .A(B0[10]), .B(w[7]), .ZN(mult_54_n703) );
  OAI22_X1 mult_54_U514 ( .A1(mult_54_n703), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n704), .ZN(mult_54_n368) );
  XNOR2_X1 mult_54_U513 ( .A(B0[9]), .B(w[7]), .ZN(mult_54_n702) );
  OAI22_X1 mult_54_U512 ( .A1(mult_54_n702), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n703), .ZN(mult_54_n369) );
  XNOR2_X1 mult_54_U511 ( .A(B0[8]), .B(w[7]), .ZN(mult_54_n701) );
  OAI22_X1 mult_54_U510 ( .A1(mult_54_n701), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n702), .ZN(mult_54_n370) );
  XNOR2_X1 mult_54_U509 ( .A(B0[7]), .B(w[7]), .ZN(mult_54_n700) );
  OAI22_X1 mult_54_U508 ( .A1(mult_54_n700), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n701), .ZN(mult_54_n371) );
  XNOR2_X1 mult_54_U507 ( .A(B0[6]), .B(w[7]), .ZN(mult_54_n699) );
  OAI22_X1 mult_54_U506 ( .A1(mult_54_n699), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n700), .ZN(mult_54_n372) );
  XNOR2_X1 mult_54_U505 ( .A(B0[5]), .B(w[7]), .ZN(mult_54_n698) );
  OAI22_X1 mult_54_U504 ( .A1(mult_54_n698), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n699), .ZN(mult_54_n373) );
  XNOR2_X1 mult_54_U503 ( .A(B0[4]), .B(w[7]), .ZN(mult_54_n697) );
  OAI22_X1 mult_54_U502 ( .A1(mult_54_n697), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n698), .ZN(mult_54_n374) );
  XNOR2_X1 mult_54_U501 ( .A(B0[3]), .B(w[7]), .ZN(mult_54_n696) );
  OAI22_X1 mult_54_U500 ( .A1(mult_54_n696), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n697), .ZN(mult_54_n375) );
  XNOR2_X1 mult_54_U499 ( .A(B0[2]), .B(w[7]), .ZN(mult_54_n695) );
  OAI22_X1 mult_54_U498 ( .A1(mult_54_n695), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n696), .ZN(mult_54_n376) );
  XNOR2_X1 mult_54_U497 ( .A(B0[1]), .B(w[7]), .ZN(mult_54_n694) );
  OAI22_X1 mult_54_U496 ( .A1(mult_54_n694), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n695), .ZN(mult_54_n377) );
  XNOR2_X1 mult_54_U495 ( .A(w[7]), .B(B0[0]), .ZN(mult_54_n692) );
  OAI22_X1 mult_54_U494 ( .A1(mult_54_n692), .A2(mult_54_n693), .B1(
        mult_54_n691), .B2(mult_54_n694), .ZN(mult_54_n378) );
  NOR2_X1 mult_54_U493 ( .A1(mult_54_n673), .A2(mult_54_n691), .ZN(
        mult_54_n379) );
  AOI21_X1 mult_54_U492 ( .B1(mult_54_n676), .B2(mult_54_n674), .A(
        mult_54_n690), .ZN(mult_54_n689) );
  INV_X1 mult_54_U491 ( .A(mult_54_n689), .ZN(mult_54_n380) );
  XNOR2_X1 mult_54_U490 ( .A(B0[11]), .B(w[5]), .ZN(mult_54_n687) );
  OAI22_X1 mult_54_U489 ( .A1(mult_54_n687), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n688), .ZN(mult_54_n381) );
  OAI22_X1 mult_54_U488 ( .A1(mult_54_n686), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n687), .ZN(mult_54_n382) );
  XNOR2_X1 mult_54_U487 ( .A(B0[8]), .B(w[5]), .ZN(mult_54_n684) );
  OAI22_X1 mult_54_U486 ( .A1(mult_54_n684), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n685), .ZN(mult_54_n384) );
  XNOR2_X1 mult_54_U485 ( .A(B0[7]), .B(w[5]), .ZN(mult_54_n683) );
  OAI22_X1 mult_54_U484 ( .A1(mult_54_n683), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n684), .ZN(mult_54_n385) );
  XNOR2_X1 mult_54_U483 ( .A(B0[6]), .B(w[5]), .ZN(mult_54_n682) );
  OAI22_X1 mult_54_U482 ( .A1(mult_54_n682), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n683), .ZN(mult_54_n386) );
  XNOR2_X1 mult_54_U481 ( .A(B0[5]), .B(w[5]), .ZN(mult_54_n681) );
  OAI22_X1 mult_54_U480 ( .A1(mult_54_n681), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n682), .ZN(mult_54_n387) );
  XNOR2_X1 mult_54_U479 ( .A(B0[4]), .B(w[5]), .ZN(mult_54_n680) );
  OAI22_X1 mult_54_U478 ( .A1(mult_54_n680), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n681), .ZN(mult_54_n388) );
  XNOR2_X1 mult_54_U477 ( .A(B0[3]), .B(w[5]), .ZN(mult_54_n679) );
  OAI22_X1 mult_54_U476 ( .A1(mult_54_n679), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n680), .ZN(mult_54_n389) );
  XNOR2_X1 mult_54_U475 ( .A(B0[2]), .B(w[5]), .ZN(mult_54_n678) );
  OAI22_X1 mult_54_U474 ( .A1(mult_54_n678), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n679), .ZN(mult_54_n390) );
  XNOR2_X1 mult_54_U473 ( .A(B0[1]), .B(w[5]), .ZN(mult_54_n677) );
  OAI22_X1 mult_54_U472 ( .A1(mult_54_n677), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n678), .ZN(mult_54_n391) );
  XNOR2_X1 mult_54_U471 ( .A(w[5]), .B(B0[0]), .ZN(mult_54_n675) );
  OAI22_X1 mult_54_U470 ( .A1(mult_54_n675), .A2(mult_54_n676), .B1(
        mult_54_n674), .B2(mult_54_n677), .ZN(mult_54_n392) );
  NOR2_X1 mult_54_U469 ( .A1(mult_54_n673), .A2(mult_54_n674), .ZN(
        mult_54_n393) );
  AOI21_X1 mult_54_U468 ( .B1(mult_54_n657), .B2(mult_54_n658), .A(
        mult_54_n672), .ZN(mult_54_n671) );
  INV_X1 mult_54_U467 ( .A(mult_54_n671), .ZN(mult_54_n394) );
  XNOR2_X1 mult_54_U466 ( .A(B0[11]), .B(w[3]), .ZN(mult_54_n669) );
  OAI22_X1 mult_54_U465 ( .A1(mult_54_n669), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n670), .ZN(mult_54_n395) );
  XNOR2_X1 mult_54_U464 ( .A(B0[10]), .B(w[3]), .ZN(mult_54_n668) );
  OAI22_X1 mult_54_U463 ( .A1(mult_54_n668), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n669), .ZN(mult_54_n396) );
  XNOR2_X1 mult_54_U462 ( .A(B0[9]), .B(w[3]), .ZN(mult_54_n667) );
  OAI22_X1 mult_54_U461 ( .A1(mult_54_n667), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n668), .ZN(mult_54_n397) );
  XNOR2_X1 mult_54_U460 ( .A(B0[8]), .B(w[3]), .ZN(mult_54_n666) );
  OAI22_X1 mult_54_U459 ( .A1(mult_54_n666), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n667), .ZN(mult_54_n398) );
  XNOR2_X1 mult_54_U458 ( .A(B0[7]), .B(w[3]), .ZN(mult_54_n665) );
  OAI22_X1 mult_54_U457 ( .A1(mult_54_n665), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n666), .ZN(mult_54_n399) );
  XNOR2_X1 mult_54_U456 ( .A(B0[6]), .B(w[3]), .ZN(mult_54_n664) );
  OAI22_X1 mult_54_U455 ( .A1(mult_54_n664), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n665), .ZN(mult_54_n400) );
  XNOR2_X1 mult_54_U454 ( .A(B0[5]), .B(w[3]), .ZN(mult_54_n663) );
  OAI22_X1 mult_54_U453 ( .A1(mult_54_n663), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n664), .ZN(mult_54_n401) );
  XNOR2_X1 mult_54_U452 ( .A(B0[4]), .B(w[3]), .ZN(mult_54_n662) );
  OAI22_X1 mult_54_U451 ( .A1(mult_54_n662), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n663), .ZN(mult_54_n402) );
  XNOR2_X1 mult_54_U450 ( .A(B0[3]), .B(w[3]), .ZN(mult_54_n661) );
  OAI22_X1 mult_54_U449 ( .A1(mult_54_n661), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n662), .ZN(mult_54_n403) );
  XNOR2_X1 mult_54_U448 ( .A(B0[2]), .B(w[3]), .ZN(mult_54_n660) );
  OAI22_X1 mult_54_U447 ( .A1(mult_54_n660), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n661), .ZN(mult_54_n404) );
  XNOR2_X1 mult_54_U446 ( .A(B0[1]), .B(w[3]), .ZN(mult_54_n659) );
  OAI22_X1 mult_54_U445 ( .A1(mult_54_n659), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n660), .ZN(mult_54_n405) );
  XNOR2_X1 mult_54_U444 ( .A(w[3]), .B(B0[0]), .ZN(mult_54_n656) );
  OAI22_X1 mult_54_U443 ( .A1(mult_54_n656), .A2(mult_54_n657), .B1(
        mult_54_n658), .B2(mult_54_n659), .ZN(mult_54_n406) );
  XOR2_X1 mult_54_U442 ( .A(B0[13]), .B(mult_54_n655), .Z(mult_54_n653) );
  AOI21_X1 mult_54_U441 ( .B1(mult_54_n641), .B2(mult_54_n643), .A(
        mult_54_n653), .ZN(mult_54_n654) );
  INV_X1 mult_54_U440 ( .A(mult_54_n654), .ZN(mult_54_n408) );
  XNOR2_X1 mult_54_U439 ( .A(B0[12]), .B(w[1]), .ZN(mult_54_n652) );
  OAI22_X1 mult_54_U438 ( .A1(mult_54_n652), .A2(mult_54_n641), .B1(
        mult_54_n653), .B2(mult_54_n643), .ZN(mult_54_n409) );
  XNOR2_X1 mult_54_U437 ( .A(B0[11]), .B(w[1]), .ZN(mult_54_n651) );
  OAI22_X1 mult_54_U436 ( .A1(mult_54_n651), .A2(mult_54_n641), .B1(
        mult_54_n652), .B2(mult_54_n643), .ZN(mult_54_n410) );
  XNOR2_X1 mult_54_U435 ( .A(B0[10]), .B(w[1]), .ZN(mult_54_n650) );
  OAI22_X1 mult_54_U434 ( .A1(mult_54_n650), .A2(mult_54_n641), .B1(
        mult_54_n651), .B2(mult_54_n643), .ZN(mult_54_n411) );
  XNOR2_X1 mult_54_U433 ( .A(B0[9]), .B(w[1]), .ZN(mult_54_n649) );
  OAI22_X1 mult_54_U432 ( .A1(mult_54_n649), .A2(mult_54_n641), .B1(
        mult_54_n650), .B2(mult_54_n643), .ZN(mult_54_n412) );
  XNOR2_X1 mult_54_U431 ( .A(B0[8]), .B(w[1]), .ZN(mult_54_n648) );
  OAI22_X1 mult_54_U430 ( .A1(mult_54_n648), .A2(mult_54_n641), .B1(
        mult_54_n649), .B2(mult_54_n643), .ZN(mult_54_n413) );
  XNOR2_X1 mult_54_U429 ( .A(B0[7]), .B(w[1]), .ZN(mult_54_n647) );
  OAI22_X1 mult_54_U428 ( .A1(mult_54_n647), .A2(mult_54_n641), .B1(
        mult_54_n648), .B2(mult_54_n643), .ZN(mult_54_n414) );
  XNOR2_X1 mult_54_U427 ( .A(B0[6]), .B(w[1]), .ZN(mult_54_n646) );
  OAI22_X1 mult_54_U426 ( .A1(mult_54_n646), .A2(mult_54_n641), .B1(
        mult_54_n647), .B2(mult_54_n643), .ZN(mult_54_n415) );
  XNOR2_X1 mult_54_U425 ( .A(B0[5]), .B(w[1]), .ZN(mult_54_n645) );
  OAI22_X1 mult_54_U424 ( .A1(mult_54_n645), .A2(mult_54_n641), .B1(
        mult_54_n646), .B2(mult_54_n643), .ZN(mult_54_n416) );
  XNOR2_X1 mult_54_U423 ( .A(B0[4]), .B(w[1]), .ZN(mult_54_n644) );
  OAI22_X1 mult_54_U422 ( .A1(mult_54_n644), .A2(mult_54_n641), .B1(
        mult_54_n645), .B2(mult_54_n643), .ZN(mult_54_n417) );
  XNOR2_X1 mult_54_U421 ( .A(B0[3]), .B(w[1]), .ZN(mult_54_n642) );
  OAI22_X1 mult_54_U420 ( .A1(mult_54_n642), .A2(mult_54_n641), .B1(
        mult_54_n644), .B2(mult_54_n643), .ZN(mult_54_n418) );
  OAI22_X1 mult_54_U419 ( .A1(mult_54_n640), .A2(mult_54_n641), .B1(
        mult_54_n642), .B2(mult_54_n643), .ZN(mult_54_n419) );
  OAI21_X1 mult_54_U418 ( .B1(mult_54_n637), .B2(mult_54_n638), .A(
        mult_54_n639), .ZN(mult_54_n636) );
  XOR2_X1 mult_54_U417 ( .A(mult_54_n636), .B(mult_54_n136), .Z(mult_54_n635)
         );
  XNOR2_X1 mult_54_U416 ( .A(mult_54_n162), .B(mult_54_n635), .ZN(temp5_26_)
         );
  XOR2_X2 mult_54_U415 ( .A(w[12]), .B(mult_54_n764), .Z(mult_54_n742) );
  XOR2_X2 mult_54_U414 ( .A(w[10]), .B(mult_54_n762), .Z(mult_54_n725) );
  XOR2_X2 mult_54_U413 ( .A(w[8]), .B(mult_54_n760), .Z(mult_54_n708) );
  XOR2_X2 mult_54_U412 ( .A(w[6]), .B(mult_54_n758), .Z(mult_54_n691) );
  XOR2_X2 mult_54_U411 ( .A(w[4]), .B(mult_54_n771), .Z(mult_54_n674) );
  INV_X1 mult_54_U410 ( .A(w[0]), .ZN(mult_54_n643) );
  INV_X1 mult_54_U409 ( .A(mult_54_n798), .ZN(mult_54_n658) );
  HA_X1 mult_54_U145 ( .A(mult_54_n406), .B(mult_54_n419), .CO(mult_54_n315), 
        .S(mult_54_n316) );
  FA_X1 mult_54_U144 ( .A(mult_54_n418), .B(mult_54_n393), .CI(mult_54_n405), 
        .CO(mult_54_n313), .S(mult_54_n314) );
  HA_X1 mult_54_U143 ( .A(mult_54_n321), .B(mult_54_n392), .CO(mult_54_n311), 
        .S(mult_54_n312) );
  FA_X1 mult_54_U142 ( .A(mult_54_n404), .B(mult_54_n417), .CI(mult_54_n312), 
        .CO(mult_54_n309), .S(mult_54_n310) );
  FA_X1 mult_54_U141 ( .A(mult_54_n416), .B(mult_54_n379), .CI(mult_54_n403), 
        .CO(mult_54_n307), .S(mult_54_n308) );
  FA_X1 mult_54_U140 ( .A(mult_54_n311), .B(mult_54_n391), .CI(mult_54_n308), 
        .CO(mult_54_n305), .S(mult_54_n306) );
  HA_X1 mult_54_U139 ( .A(mult_54_n320), .B(mult_54_n378), .CO(mult_54_n303), 
        .S(mult_54_n304) );
  FA_X1 mult_54_U138 ( .A(mult_54_n390), .B(mult_54_n415), .CI(mult_54_n402), 
        .CO(mult_54_n301), .S(mult_54_n302) );
  FA_X1 mult_54_U137 ( .A(mult_54_n307), .B(mult_54_n304), .CI(mult_54_n302), 
        .CO(mult_54_n299), .S(mult_54_n300) );
  FA_X1 mult_54_U136 ( .A(mult_54_n389), .B(mult_54_n365), .CI(mult_54_n414), 
        .CO(mult_54_n297), .S(mult_54_n298) );
  FA_X1 mult_54_U135 ( .A(mult_54_n377), .B(mult_54_n401), .CI(mult_54_n303), 
        .CO(mult_54_n295), .S(mult_54_n296) );
  FA_X1 mult_54_U134 ( .A(mult_54_n298), .B(mult_54_n301), .CI(mult_54_n296), 
        .CO(mult_54_n293), .S(mult_54_n294) );
  HA_X1 mult_54_U133 ( .A(mult_54_n319), .B(mult_54_n364), .CO(mult_54_n291), 
        .S(mult_54_n292) );
  FA_X1 mult_54_U132 ( .A(mult_54_n376), .B(mult_54_n388), .CI(mult_54_n400), 
        .CO(mult_54_n289), .S(mult_54_n290) );
  FA_X1 mult_54_U131 ( .A(mult_54_n292), .B(mult_54_n413), .CI(mult_54_n297), 
        .CO(mult_54_n287), .S(mult_54_n288) );
  FA_X1 mult_54_U130 ( .A(mult_54_n290), .B(mult_54_n295), .CI(mult_54_n288), 
        .CO(mult_54_n285), .S(mult_54_n286) );
  FA_X1 mult_54_U129 ( .A(mult_54_n375), .B(mult_54_n351), .CI(mult_54_n412), 
        .CO(mult_54_n283), .S(mult_54_n284) );
  FA_X1 mult_54_U128 ( .A(mult_54_n363), .B(mult_54_n399), .CI(mult_54_n387), 
        .CO(mult_54_n281), .S(mult_54_n282) );
  FA_X1 mult_54_U127 ( .A(mult_54_n289), .B(mult_54_n291), .CI(mult_54_n284), 
        .CO(mult_54_n279), .S(mult_54_n280) );
  FA_X1 mult_54_U126 ( .A(mult_54_n287), .B(mult_54_n282), .CI(mult_54_n280), 
        .CO(mult_54_n277), .S(mult_54_n278) );
  HA_X1 mult_54_U125 ( .A(mult_54_n318), .B(mult_54_n350), .CO(mult_54_n275), 
        .S(mult_54_n276) );
  FA_X1 mult_54_U124 ( .A(mult_54_n362), .B(mult_54_n386), .CI(mult_54_n411), 
        .CO(mult_54_n273), .S(mult_54_n274) );
  FA_X1 mult_54_U123 ( .A(mult_54_n374), .B(mult_54_n398), .CI(mult_54_n276), 
        .CO(mult_54_n271), .S(mult_54_n272) );
  FA_X1 mult_54_U122 ( .A(mult_54_n281), .B(mult_54_n283), .CI(mult_54_n274), 
        .CO(mult_54_n269), .S(mult_54_n270) );
  FA_X1 mult_54_U121 ( .A(mult_54_n279), .B(mult_54_n272), .CI(mult_54_n270), 
        .CO(mult_54_n267), .S(mult_54_n268) );
  FA_X1 mult_54_U120 ( .A(mult_54_n361), .B(mult_54_n337), .CI(mult_54_n410), 
        .CO(mult_54_n265), .S(mult_54_n266) );
  FA_X1 mult_54_U109 ( .A(mult_54_n349), .B(mult_54_n397), .CI(mult_54_n373), 
        .CO(mult_54_n263), .S(mult_54_n264) );
  FA_X1 mult_54_U108 ( .A(mult_54_n275), .B(mult_54_n385), .CI(mult_54_n273), 
        .CO(mult_54_n261), .S(mult_54_n262) );
  FA_X1 mult_54_U107 ( .A(mult_54_n264), .B(mult_54_n266), .CI(mult_54_n271), 
        .CO(mult_54_n259), .S(mult_54_n260) );
  FA_X1 mult_54_U106 ( .A(mult_54_n262), .B(mult_54_n269), .CI(mult_54_n260), 
        .CO(mult_54_n257), .S(mult_54_n258) );
  HA_X1 mult_54_U105 ( .A(mult_54_n317), .B(mult_54_n336), .CO(mult_54_n255), 
        .S(mult_54_n256) );
  FA_X1 mult_54_U104 ( .A(mult_54_n409), .B(mult_54_n372), .CI(mult_54_n396), 
        .CO(mult_54_n253), .S(mult_54_n254) );
  FA_X1 mult_54_U103 ( .A(mult_54_n348), .B(mult_54_n384), .CI(mult_54_n360), 
        .CO(mult_54_n251), .S(mult_54_n252) );
  FA_X1 mult_54_U102 ( .A(mult_54_n265), .B(mult_54_n256), .CI(mult_54_n263), 
        .CO(mult_54_n249), .S(mult_54_n250) );
  FA_X1 mult_54_U101 ( .A(mult_54_n254), .B(mult_54_n252), .CI(mult_54_n261), 
        .CO(mult_54_n247), .S(mult_54_n248) );
  FA_X1 mult_54_U100 ( .A(mult_54_n259), .B(mult_54_n250), .CI(mult_54_n248), 
        .CO(mult_54_n245), .S(mult_54_n246) );
  FA_X1 mult_54_U97 ( .A(mult_54_n395), .B(mult_54_n359), .CI(mult_54_n408), 
        .CO(mult_54_n241), .S(mult_54_n242) );
  FA_X1 mult_54_U96 ( .A(mult_54_n335), .B(mult_54_n371), .CI(mult_54_n255), 
        .CO(mult_54_n239), .S(mult_54_n240) );
  FA_X1 mult_54_U95 ( .A(mult_54_n253), .B(mult_54_n244), .CI(mult_54_n251), 
        .CO(mult_54_n237), .S(mult_54_n238) );
  FA_X1 mult_54_U94 ( .A(mult_54_n240), .B(mult_54_n242), .CI(mult_54_n249), 
        .CO(mult_54_n235), .S(mult_54_n236) );
  FA_X1 mult_54_U93 ( .A(mult_54_n247), .B(mult_54_n238), .CI(mult_54_n236), 
        .CO(mult_54_n233), .S(mult_54_n234) );
  FA_X1 mult_54_U91 ( .A(mult_54_n382), .B(mult_54_n346), .CI(mult_54_n232), 
        .CO(mult_54_n229), .S(mult_54_n230) );
  FA_X1 mult_54_U90 ( .A(mult_54_n334), .B(mult_54_n370), .CI(mult_54_n358), 
        .CO(mult_54_n227), .S(mult_54_n228) );
  FA_X1 mult_54_U89 ( .A(mult_54_n241), .B(mult_54_n243), .CI(mult_54_n239), 
        .CO(mult_54_n225), .S(mult_54_n226) );
  FA_X1 mult_54_U88 ( .A(mult_54_n230), .B(mult_54_n228), .CI(mult_54_n237), 
        .CO(mult_54_n223), .S(mult_54_n224) );
  FA_X1 mult_54_U87 ( .A(mult_54_n235), .B(mult_54_n226), .CI(mult_54_n224), 
        .CO(mult_54_n221), .S(mult_54_n222) );
  FA_X1 mult_54_U86 ( .A(mult_54_n231), .B(mult_54_n333), .CI(mult_54_n394), 
        .CO(mult_54_n219), .S(mult_54_n220) );
  FA_X1 mult_54_U85 ( .A(mult_54_n345), .B(mult_54_n381), .CI(mult_54_n357), 
        .CO(mult_54_n217), .S(mult_54_n218) );
  FA_X1 mult_54_U84 ( .A(mult_54_n229), .B(mult_54_n369), .CI(mult_54_n227), 
        .CO(mult_54_n215), .S(mult_54_n216) );
  FA_X1 mult_54_U83 ( .A(mult_54_n220), .B(mult_54_n218), .CI(mult_54_n225), 
        .CO(mult_54_n213), .S(mult_54_n214) );
  FA_X1 mult_54_U82 ( .A(mult_54_n223), .B(mult_54_n216), .CI(mult_54_n214), 
        .CO(mult_54_n211), .S(mult_54_n212) );
  FA_X1 mult_54_U80 ( .A(mult_54_n368), .B(mult_54_n344), .CI(mult_54_n210), 
        .CO(mult_54_n207), .S(mult_54_n208) );
  FA_X1 mult_54_U79 ( .A(mult_54_n332), .B(mult_54_n356), .CI(mult_54_n219), 
        .CO(mult_54_n205), .S(mult_54_n206) );
  FA_X1 mult_54_U78 ( .A(mult_54_n208), .B(mult_54_n217), .CI(mult_54_n215), 
        .CO(mult_54_n203), .S(mult_54_n204) );
  FA_X1 mult_54_U77 ( .A(mult_54_n213), .B(mult_54_n206), .CI(mult_54_n204), 
        .CO(mult_54_n201), .S(mult_54_n202) );
  FA_X1 mult_54_U76 ( .A(mult_54_n209), .B(mult_54_n331), .CI(mult_54_n380), 
        .CO(mult_54_n199), .S(mult_54_n200) );
  FA_X1 mult_54_U75 ( .A(mult_54_n355), .B(mult_54_n343), .CI(mult_54_n367), 
        .CO(mult_54_n197), .S(mult_54_n198) );
  FA_X1 mult_54_U74 ( .A(mult_54_n198), .B(mult_54_n207), .CI(mult_54_n200), 
        .CO(mult_54_n195), .S(mult_54_n196) );
  FA_X1 mult_54_U73 ( .A(mult_54_n203), .B(mult_54_n205), .CI(mult_54_n196), 
        .CO(mult_54_n193), .S(mult_54_n194) );
  FA_X1 mult_54_U71 ( .A(mult_54_n330), .B(mult_54_n342), .CI(mult_54_n192), 
        .CO(mult_54_n189), .S(mult_54_n190) );
  FA_X1 mult_54_U70 ( .A(mult_54_n199), .B(mult_54_n354), .CI(mult_54_n197), 
        .CO(mult_54_n187), .S(mult_54_n188) );
  FA_X1 mult_54_U69 ( .A(mult_54_n188), .B(mult_54_n190), .CI(mult_54_n195), 
        .CO(mult_54_n185), .S(mult_54_n186) );
  FA_X1 mult_54_U68 ( .A(mult_54_n191), .B(mult_54_n329), .CI(mult_54_n366), 
        .CO(mult_54_n183), .S(mult_54_n184) );
  FA_X1 mult_54_U67 ( .A(mult_54_n341), .B(mult_54_n353), .CI(mult_54_n189), 
        .CO(mult_54_n181), .S(mult_54_n182) );
  FA_X1 mult_54_U66 ( .A(mult_54_n187), .B(mult_54_n184), .CI(mult_54_n182), 
        .CO(mult_54_n179), .S(mult_54_n180) );
  FA_X1 mult_54_U64 ( .A(mult_54_n328), .B(mult_54_n340), .CI(mult_54_n178), 
        .CO(mult_54_n175), .S(mult_54_n176) );
  FA_X1 mult_54_U63 ( .A(mult_54_n176), .B(mult_54_n183), .CI(mult_54_n181), 
        .CO(mult_54_n173), .S(mult_54_n174) );
  FA_X1 mult_54_U62 ( .A(mult_54_n327), .B(mult_54_n177), .CI(mult_54_n352), 
        .CO(mult_54_n171), .S(mult_54_n172) );
  FA_X1 mult_54_U61 ( .A(mult_54_n175), .B(mult_54_n339), .CI(mult_54_n172), 
        .CO(mult_54_n169), .S(mult_54_n170) );
  FA_X1 mult_54_U59 ( .A(mult_54_n168), .B(mult_54_n326), .CI(mult_54_n171), 
        .CO(mult_54_n165), .S(mult_54_n166) );
  FA_X1 mult_54_U58 ( .A(mult_54_n325), .B(mult_54_n167), .CI(mult_54_n338), 
        .CO(mult_54_n163), .S(mult_54_n164) );
  FA_X1 mult_54_U44 ( .A(mult_54_n246), .B(mult_54_n257), .CI(mult_54_n149), 
        .CO(mult_54_n148), .S(temp5_13_) );
  FA_X1 mult_54_U43 ( .A(mult_54_n234), .B(mult_54_n245), .CI(mult_54_n148), 
        .CO(mult_54_n147), .S(temp5_14_) );
  FA_X1 mult_54_U42 ( .A(mult_54_n222), .B(mult_54_n233), .CI(mult_54_n147), 
        .CO(mult_54_n146), .S(temp5_15_) );
  FA_X1 mult_54_U41 ( .A(mult_54_n212), .B(mult_54_n221), .CI(mult_54_n146), 
        .CO(mult_54_n145), .S(temp5_16_) );
  FA_X1 mult_54_U40 ( .A(mult_54_n202), .B(mult_54_n211), .CI(mult_54_n145), 
        .CO(mult_54_n144), .S(temp5_17_) );
  FA_X1 mult_54_U39 ( .A(mult_54_n194), .B(mult_54_n201), .CI(mult_54_n144), 
        .CO(mult_54_n143), .S(temp5_18_) );
  FA_X1 mult_54_U38 ( .A(mult_54_n186), .B(mult_54_n193), .CI(mult_54_n143), 
        .CO(mult_54_n142), .S(temp5_19_) );
  FA_X1 mult_54_U37 ( .A(mult_54_n180), .B(mult_54_n185), .CI(mult_54_n142), 
        .CO(mult_54_n141), .S(temp5_20_) );
  FA_X1 mult_54_U30 ( .A(mult_54_n174), .B(mult_54_n179), .CI(mult_54_n141), 
        .CO(mult_54_n140), .S(temp5_21_) );
  FA_X1 mult_54_U20 ( .A(mult_54_n170), .B(mult_54_n173), .CI(mult_54_n140), 
        .CO(mult_54_n139), .S(temp5_22_) );
  FA_X1 mult_54_U10 ( .A(mult_54_n166), .B(mult_54_n169), .CI(mult_54_n139), 
        .CO(mult_54_n138), .S(temp5_23_) );
  FA_X1 mult_54_U9 ( .A(mult_54_n165), .B(mult_54_n164), .CI(mult_54_n138), 
        .CO(mult_54_n137), .S(temp5_24_) );
  FA_X1 mult_54_U8 ( .A(mult_54_n163), .B(mult_54_n162), .CI(mult_54_n137), 
        .CO(mult_54_n136), .S(temp5_25_) );
  XOR2_X1 add_0_root_add_0_root_add_59_U2 ( .A(temp5_13_), .B(ff_0_), .Z(
        DOUT[0]) );
  AND2_X1 add_0_root_add_0_root_add_59_U1 ( .A1(ff_0_), .A2(temp5_13_), .ZN(
        add_0_root_add_0_root_add_59_carry_1_) );
  FA_X1 add_0_root_add_0_root_add_59_U1_1 ( .A(ff_1_), .B(temp5_14_), .CI(
        add_0_root_add_0_root_add_59_carry_1_), .CO(
        add_0_root_add_0_root_add_59_carry_2_), .S(DOUT[1]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_2 ( .A(ff_2_), .B(temp5_15_), .CI(
        add_0_root_add_0_root_add_59_carry_2_), .CO(
        add_0_root_add_0_root_add_59_carry_3_), .S(DOUT[2]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_3 ( .A(ff_3_), .B(temp5_16_), .CI(
        add_0_root_add_0_root_add_59_carry_3_), .CO(
        add_0_root_add_0_root_add_59_carry_4_), .S(DOUT[3]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_4 ( .A(ff_4_), .B(temp5_17_), .CI(
        add_0_root_add_0_root_add_59_carry_4_), .CO(
        add_0_root_add_0_root_add_59_carry_5_), .S(DOUT[4]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_5 ( .A(ff_5_), .B(temp5_18_), .CI(
        add_0_root_add_0_root_add_59_carry_5_), .CO(
        add_0_root_add_0_root_add_59_carry_6_), .S(DOUT[5]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_6 ( .A(ff_6_), .B(temp5_19_), .CI(
        add_0_root_add_0_root_add_59_carry_6_), .CO(
        add_0_root_add_0_root_add_59_carry_7_), .S(DOUT[6]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_7 ( .A(ff_7_), .B(temp5_20_), .CI(
        add_0_root_add_0_root_add_59_carry_7_), .CO(
        add_0_root_add_0_root_add_59_carry_8_), .S(DOUT[7]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_8 ( .A(ff_8_), .B(temp5_21_), .CI(
        add_0_root_add_0_root_add_59_carry_8_), .CO(
        add_0_root_add_0_root_add_59_carry_9_), .S(DOUT[8]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_9 ( .A(ff_9_), .B(temp5_22_), .CI(
        add_0_root_add_0_root_add_59_carry_9_), .CO(
        add_0_root_add_0_root_add_59_carry_10_), .S(DOUT[9]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_10 ( .A(ff_10_), .B(temp5_23_), .CI(
        add_0_root_add_0_root_add_59_carry_10_), .CO(
        add_0_root_add_0_root_add_59_carry_11_), .S(DOUT[10]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_11 ( .A(ff_11_), .B(temp5_24_), .CI(
        add_0_root_add_0_root_add_59_carry_11_), .CO(
        add_0_root_add_0_root_add_59_carry_12_), .S(DOUT[11]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_12 ( .A(ff_12_), .B(temp5_25_), .CI(
        add_0_root_add_0_root_add_59_carry_12_), .CO(
        add_0_root_add_0_root_add_59_carry_13_), .S(DOUT[12]) );
  FA_X1 add_0_root_add_0_root_add_59_U1_13 ( .A(ff_13_), .B(temp5_26_), .CI(
        add_0_root_add_0_root_add_59_carry_13_), .S(DOUT[13]) );
  XOR2_X1 mult_46_U698 ( .A(reg1[2]), .B(mult_46_n635), .Z(mult_46_n805) );
  NOR2_X1 mult_46_U697 ( .A1(mult_46_n636), .A2(A1[1]), .ZN(mult_46_n810) );
  INV_X1 mult_46_U696 ( .A(mult_46_n810), .ZN(mult_46_n812) );
  NAND2_X1 mult_46_U695 ( .A1(n172), .A2(mult_46_n657), .ZN(mult_46_n655) );
  XNOR2_X1 mult_46_U694 ( .A(A1[2]), .B(mult_46_n635), .ZN(mult_46_n654) );
  OAI22_X1 mult_46_U693 ( .A1(mult_46_n812), .A2(mult_46_n655), .B1(
        mult_46_n654), .B2(mult_46_n657), .ZN(mult_46_n811) );
  NAND2_X1 mult_46_U692 ( .A1(mult_46_n805), .A2(mult_46_n811), .ZN(
        mult_46_n808) );
  NAND2_X1 mult_46_U691 ( .A1(mult_46_n810), .A2(mult_46_n811), .ZN(
        mult_46_n809) );
  INV_X1 mult_46_U690 ( .A(A1[0]), .ZN(mult_46_n686) );
  MUX2_X1 mult_46_U689 ( .A(mult_46_n808), .B(mult_46_n809), .S(mult_46_n686), 
        .Z(mult_46_n807) );
  INV_X1 mult_46_U688 ( .A(mult_46_n807), .ZN(mult_46_n802) );
  XNOR2_X1 mult_46_U687 ( .A(mult_46_n638), .B(reg1[2]), .ZN(mult_46_n806) );
  NAND2_X1 mult_46_U686 ( .A1(mult_46_n671), .A2(mult_46_n806), .ZN(
        mult_46_n670) );
  NAND3_X1 mult_46_U685 ( .A1(mult_46_n805), .A2(mult_46_n686), .A3(
        mult_46_n637), .ZN(mult_46_n804) );
  OAI21_X1 mult_46_U684 ( .B1(mult_46_n638), .B2(mult_46_n670), .A(
        mult_46_n804), .ZN(mult_46_n803) );
  AOI222_X1 mult_46_U683 ( .A1(mult_46_n802), .A2(mult_46_n316), .B1(
        mult_46_n803), .B2(mult_46_n802), .C1(mult_46_n803), .C2(mult_46_n316), 
        .ZN(mult_46_n801) );
  INV_X1 mult_46_U682 ( .A(mult_46_n801), .ZN(mult_46_n800) );
  AOI222_X1 mult_46_U681 ( .A1(mult_46_n800), .A2(mult_46_n314), .B1(
        mult_46_n800), .B2(mult_46_n315), .C1(mult_46_n315), .C2(mult_46_n314), 
        .ZN(mult_46_n799) );
  INV_X1 mult_46_U680 ( .A(mult_46_n799), .ZN(mult_46_n798) );
  AOI222_X1 mult_46_U679 ( .A1(mult_46_n798), .A2(mult_46_n310), .B1(
        mult_46_n798), .B2(mult_46_n313), .C1(mult_46_n313), .C2(mult_46_n310), 
        .ZN(mult_46_n797) );
  INV_X1 mult_46_U678 ( .A(mult_46_n797), .ZN(mult_46_n796) );
  AOI222_X1 mult_46_U677 ( .A1(mult_46_n796), .A2(mult_46_n306), .B1(
        mult_46_n796), .B2(mult_46_n309), .C1(mult_46_n309), .C2(mult_46_n306), 
        .ZN(mult_46_n795) );
  INV_X1 mult_46_U676 ( .A(mult_46_n795), .ZN(mult_46_n794) );
  AOI222_X1 mult_46_U675 ( .A1(mult_46_n794), .A2(mult_46_n300), .B1(
        mult_46_n794), .B2(mult_46_n305), .C1(mult_46_n305), .C2(mult_46_n300), 
        .ZN(mult_46_n793) );
  INV_X1 mult_46_U674 ( .A(mult_46_n793), .ZN(mult_46_n792) );
  AOI222_X1 mult_46_U673 ( .A1(mult_46_n792), .A2(mult_46_n294), .B1(
        mult_46_n792), .B2(mult_46_n299), .C1(mult_46_n299), .C2(mult_46_n294), 
        .ZN(mult_46_n791) );
  INV_X1 mult_46_U672 ( .A(mult_46_n791), .ZN(mult_46_n790) );
  AOI222_X1 mult_46_U671 ( .A1(mult_46_n790), .A2(mult_46_n286), .B1(
        mult_46_n790), .B2(mult_46_n293), .C1(mult_46_n293), .C2(mult_46_n286), 
        .ZN(mult_46_n787) );
  INV_X1 mult_46_U670 ( .A(mult_46_n278), .ZN(mult_46_n788) );
  INV_X1 mult_46_U669 ( .A(mult_46_n285), .ZN(mult_46_n789) );
  OAI222_X1 mult_46_U668 ( .A1(mult_46_n787), .A2(mult_46_n788), .B1(
        mult_46_n787), .B2(mult_46_n789), .C1(mult_46_n789), .C2(mult_46_n788), 
        .ZN(mult_46_n786) );
  AOI222_X1 mult_46_U667 ( .A1(mult_46_n786), .A2(mult_46_n268), .B1(
        mult_46_n786), .B2(mult_46_n277), .C1(mult_46_n277), .C2(mult_46_n268), 
        .ZN(mult_46_n783) );
  INV_X1 mult_46_U666 ( .A(mult_46_n258), .ZN(mult_46_n784) );
  INV_X1 mult_46_U665 ( .A(mult_46_n267), .ZN(mult_46_n785) );
  OAI222_X1 mult_46_U664 ( .A1(mult_46_n783), .A2(mult_46_n784), .B1(
        mult_46_n783), .B2(mult_46_n785), .C1(mult_46_n785), .C2(mult_46_n784), 
        .ZN(mult_46_n149) );
  XOR2_X1 mult_46_U663 ( .A(A1[12]), .B(mult_46_n647), .Z(mult_46_n770) );
  XNOR2_X1 mult_46_U662 ( .A(mult_46_n648), .B(reg1[12]), .ZN(mult_46_n782) );
  NAND2_X1 mult_46_U661 ( .A1(mult_46_n755), .A2(mult_46_n782), .ZN(
        mult_46_n757) );
  INV_X1 mult_46_U660 ( .A(mult_46_n757), .ZN(mult_46_n651) );
  INV_X1 mult_46_U659 ( .A(mult_46_n755), .ZN(mult_46_n652) );
  XNOR2_X1 mult_46_U658 ( .A(A1[13]), .B(mult_46_n648), .ZN(mult_46_n653) );
  AOI22_X1 mult_46_U657 ( .A1(mult_46_n770), .A2(mult_46_n651), .B1(
        mult_46_n652), .B2(mult_46_n653), .ZN(mult_46_n162) );
  XNOR2_X1 mult_46_U656 ( .A(A1[12]), .B(mult_46_n645), .ZN(mult_46_n752) );
  XNOR2_X1 mult_46_U655 ( .A(mult_46_n646), .B(reg1[10]), .ZN(mult_46_n781) );
  NAND2_X1 mult_46_U654 ( .A1(mult_46_n738), .A2(mult_46_n781), .ZN(
        mult_46_n740) );
  XNOR2_X1 mult_46_U653 ( .A(A1[13]), .B(mult_46_n645), .ZN(mult_46_n754) );
  OAI22_X1 mult_46_U652 ( .A1(mult_46_n752), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n754), .ZN(mult_46_n167) );
  INV_X1 mult_46_U651 ( .A(mult_46_n167), .ZN(mult_46_n168) );
  XNOR2_X1 mult_46_U650 ( .A(A1[12]), .B(mult_46_n643), .ZN(mult_46_n735) );
  XNOR2_X1 mult_46_U649 ( .A(mult_46_n644), .B(reg1[8]), .ZN(mult_46_n780) );
  NAND2_X1 mult_46_U648 ( .A1(mult_46_n721), .A2(mult_46_n780), .ZN(
        mult_46_n723) );
  XNOR2_X1 mult_46_U647 ( .A(A1[13]), .B(mult_46_n643), .ZN(mult_46_n737) );
  OAI22_X1 mult_46_U646 ( .A1(mult_46_n735), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n737), .ZN(mult_46_n177) );
  INV_X1 mult_46_U645 ( .A(mult_46_n177), .ZN(mult_46_n178) );
  XNOR2_X1 mult_46_U644 ( .A(A1[12]), .B(mult_46_n641), .ZN(mult_46_n718) );
  XNOR2_X1 mult_46_U643 ( .A(mult_46_n642), .B(reg1[6]), .ZN(mult_46_n779) );
  NAND2_X1 mult_46_U642 ( .A1(mult_46_n704), .A2(mult_46_n779), .ZN(
        mult_46_n706) );
  XNOR2_X1 mult_46_U641 ( .A(A1[13]), .B(mult_46_n641), .ZN(mult_46_n720) );
  OAI22_X1 mult_46_U640 ( .A1(mult_46_n718), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n720), .ZN(mult_46_n191) );
  INV_X1 mult_46_U639 ( .A(mult_46_n191), .ZN(mult_46_n192) );
  XNOR2_X1 mult_46_U638 ( .A(A1[12]), .B(mult_46_n639), .ZN(mult_46_n701) );
  XNOR2_X1 mult_46_U637 ( .A(mult_46_n640), .B(reg1[4]), .ZN(mult_46_n778) );
  NAND2_X1 mult_46_U636 ( .A1(mult_46_n687), .A2(mult_46_n778), .ZN(
        mult_46_n689) );
  XNOR2_X1 mult_46_U635 ( .A(A1[13]), .B(mult_46_n639), .ZN(mult_46_n703) );
  OAI22_X1 mult_46_U634 ( .A1(mult_46_n701), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n703), .ZN(mult_46_n209) );
  INV_X1 mult_46_U633 ( .A(mult_46_n209), .ZN(mult_46_n210) );
  XNOR2_X1 mult_46_U632 ( .A(A1[12]), .B(mult_46_n637), .ZN(mult_46_n683) );
  XNOR2_X1 mult_46_U631 ( .A(A1[13]), .B(mult_46_n637), .ZN(mult_46_n685) );
  OAI22_X1 mult_46_U630 ( .A1(mult_46_n683), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n685), .ZN(mult_46_n231) );
  INV_X1 mult_46_U629 ( .A(mult_46_n231), .ZN(mult_46_n232) );
  XNOR2_X1 mult_46_U628 ( .A(A1[3]), .B(mult_46_n645), .ZN(mult_46_n743) );
  XNOR2_X1 mult_46_U627 ( .A(A1[4]), .B(mult_46_n645), .ZN(mult_46_n744) );
  OAI22_X1 mult_46_U626 ( .A1(mult_46_n743), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n744), .ZN(mult_46_n776) );
  XNOR2_X1 mult_46_U625 ( .A(A1[9]), .B(mult_46_n639), .ZN(mult_46_n698) );
  XNOR2_X1 mult_46_U624 ( .A(A1[10]), .B(mult_46_n639), .ZN(mult_46_n699) );
  OAI22_X1 mult_46_U623 ( .A1(mult_46_n698), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n699), .ZN(mult_46_n777) );
  OR2_X1 mult_46_U622 ( .A1(mult_46_n776), .A2(mult_46_n777), .ZN(mult_46_n243) );
  XNOR2_X1 mult_46_U621 ( .A(mult_46_n776), .B(mult_46_n777), .ZN(mult_46_n244) );
  NAND3_X1 mult_46_U620 ( .A1(mult_46_n652), .A2(mult_46_n686), .A3(n184), 
        .ZN(mult_46_n775) );
  OAI21_X1 mult_46_U619 ( .B1(mult_46_n648), .B2(mult_46_n757), .A(
        mult_46_n775), .ZN(mult_46_n317) );
  OR3_X1 mult_46_U618 ( .A1(mult_46_n738), .A2(A1[0]), .A3(mult_46_n646), .ZN(
        mult_46_n774) );
  OAI21_X1 mult_46_U617 ( .B1(mult_46_n646), .B2(mult_46_n740), .A(
        mult_46_n774), .ZN(mult_46_n318) );
  OR3_X1 mult_46_U616 ( .A1(mult_46_n721), .A2(A1[0]), .A3(mult_46_n644), .ZN(
        mult_46_n773) );
  OAI21_X1 mult_46_U615 ( .B1(mult_46_n644), .B2(mult_46_n723), .A(
        mult_46_n773), .ZN(mult_46_n319) );
  OR3_X1 mult_46_U614 ( .A1(mult_46_n704), .A2(A1[0]), .A3(mult_46_n642), .ZN(
        mult_46_n772) );
  OAI21_X1 mult_46_U613 ( .B1(mult_46_n642), .B2(mult_46_n706), .A(
        mult_46_n772), .ZN(mult_46_n320) );
  OR3_X1 mult_46_U612 ( .A1(mult_46_n687), .A2(A1[0]), .A3(mult_46_n640), .ZN(
        mult_46_n771) );
  OAI21_X1 mult_46_U611 ( .B1(mult_46_n640), .B2(mult_46_n689), .A(
        mult_46_n771), .ZN(mult_46_n321) );
  XNOR2_X1 mult_46_U610 ( .A(A1[11]), .B(mult_46_n647), .ZN(mult_46_n768) );
  INV_X1 mult_46_U609 ( .A(mult_46_n770), .ZN(mult_46_n769) );
  OAI22_X1 mult_46_U608 ( .A1(mult_46_n768), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n769), .ZN(mult_46_n325) );
  XNOR2_X1 mult_46_U607 ( .A(A1[10]), .B(mult_46_n647), .ZN(mult_46_n767) );
  OAI22_X1 mult_46_U606 ( .A1(mult_46_n767), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n768), .ZN(mult_46_n326) );
  XNOR2_X1 mult_46_U605 ( .A(A1[9]), .B(mult_46_n647), .ZN(mult_46_n766) );
  OAI22_X1 mult_46_U604 ( .A1(mult_46_n766), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n767), .ZN(mult_46_n327) );
  XNOR2_X1 mult_46_U603 ( .A(A1[8]), .B(mult_46_n647), .ZN(mult_46_n765) );
  OAI22_X1 mult_46_U602 ( .A1(mult_46_n765), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n766), .ZN(mult_46_n328) );
  XNOR2_X1 mult_46_U601 ( .A(A1[7]), .B(mult_46_n647), .ZN(mult_46_n764) );
  OAI22_X1 mult_46_U600 ( .A1(mult_46_n764), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n765), .ZN(mult_46_n329) );
  XNOR2_X1 mult_46_U599 ( .A(A1[6]), .B(mult_46_n647), .ZN(mult_46_n763) );
  OAI22_X1 mult_46_U598 ( .A1(mult_46_n763), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n764), .ZN(mult_46_n330) );
  XNOR2_X1 mult_46_U597 ( .A(A1[5]), .B(mult_46_n647), .ZN(mult_46_n762) );
  OAI22_X1 mult_46_U596 ( .A1(mult_46_n762), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n763), .ZN(mult_46_n331) );
  XNOR2_X1 mult_46_U595 ( .A(A1[4]), .B(mult_46_n647), .ZN(mult_46_n761) );
  OAI22_X1 mult_46_U594 ( .A1(mult_46_n761), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n762), .ZN(mult_46_n332) );
  XNOR2_X1 mult_46_U593 ( .A(A1[3]), .B(mult_46_n647), .ZN(mult_46_n760) );
  OAI22_X1 mult_46_U592 ( .A1(mult_46_n760), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n761), .ZN(mult_46_n333) );
  XNOR2_X1 mult_46_U591 ( .A(A1[2]), .B(mult_46_n647), .ZN(mult_46_n759) );
  OAI22_X1 mult_46_U590 ( .A1(mult_46_n759), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n760), .ZN(mult_46_n334) );
  XNOR2_X1 mult_46_U589 ( .A(A1[1]), .B(mult_46_n647), .ZN(mult_46_n758) );
  OAI22_X1 mult_46_U588 ( .A1(mult_46_n758), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n759), .ZN(mult_46_n335) );
  XNOR2_X1 mult_46_U587 ( .A(n184), .B(A1[0]), .ZN(mult_46_n756) );
  OAI22_X1 mult_46_U586 ( .A1(mult_46_n756), .A2(mult_46_n757), .B1(
        mult_46_n755), .B2(mult_46_n758), .ZN(mult_46_n336) );
  NOR2_X1 mult_46_U585 ( .A1(mult_46_n686), .A2(mult_46_n755), .ZN(
        mult_46_n337) );
  AOI21_X1 mult_46_U584 ( .B1(mult_46_n740), .B2(mult_46_n738), .A(
        mult_46_n754), .ZN(mult_46_n753) );
  INV_X1 mult_46_U583 ( .A(mult_46_n753), .ZN(mult_46_n338) );
  XNOR2_X1 mult_46_U582 ( .A(A1[11]), .B(mult_46_n645), .ZN(mult_46_n751) );
  OAI22_X1 mult_46_U581 ( .A1(mult_46_n751), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n752), .ZN(mult_46_n339) );
  XNOR2_X1 mult_46_U580 ( .A(A1[10]), .B(mult_46_n645), .ZN(mult_46_n750) );
  OAI22_X1 mult_46_U579 ( .A1(mult_46_n750), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n751), .ZN(mult_46_n340) );
  XNOR2_X1 mult_46_U578 ( .A(A1[9]), .B(mult_46_n645), .ZN(mult_46_n749) );
  OAI22_X1 mult_46_U577 ( .A1(mult_46_n749), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n750), .ZN(mult_46_n341) );
  XNOR2_X1 mult_46_U576 ( .A(A1[8]), .B(mult_46_n645), .ZN(mult_46_n748) );
  OAI22_X1 mult_46_U575 ( .A1(mult_46_n748), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n749), .ZN(mult_46_n342) );
  XNOR2_X1 mult_46_U574 ( .A(A1[7]), .B(mult_46_n645), .ZN(mult_46_n747) );
  OAI22_X1 mult_46_U573 ( .A1(mult_46_n747), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n748), .ZN(mult_46_n343) );
  XNOR2_X1 mult_46_U572 ( .A(A1[6]), .B(mult_46_n645), .ZN(mult_46_n746) );
  OAI22_X1 mult_46_U571 ( .A1(mult_46_n746), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n747), .ZN(mult_46_n344) );
  XNOR2_X1 mult_46_U570 ( .A(A1[5]), .B(mult_46_n645), .ZN(mult_46_n745) );
  OAI22_X1 mult_46_U569 ( .A1(mult_46_n745), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n746), .ZN(mult_46_n345) );
  OAI22_X1 mult_46_U568 ( .A1(mult_46_n744), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n745), .ZN(mult_46_n346) );
  XNOR2_X1 mult_46_U567 ( .A(A1[2]), .B(mult_46_n645), .ZN(mult_46_n742) );
  OAI22_X1 mult_46_U566 ( .A1(mult_46_n742), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n743), .ZN(mult_46_n348) );
  XNOR2_X1 mult_46_U565 ( .A(A1[1]), .B(mult_46_n645), .ZN(mult_46_n741) );
  OAI22_X1 mult_46_U564 ( .A1(mult_46_n741), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n742), .ZN(mult_46_n349) );
  XNOR2_X1 mult_46_U563 ( .A(n182), .B(A1[0]), .ZN(mult_46_n739) );
  OAI22_X1 mult_46_U562 ( .A1(mult_46_n739), .A2(mult_46_n740), .B1(
        mult_46_n738), .B2(mult_46_n741), .ZN(mult_46_n350) );
  NOR2_X1 mult_46_U561 ( .A1(mult_46_n686), .A2(mult_46_n738), .ZN(
        mult_46_n351) );
  AOI21_X1 mult_46_U560 ( .B1(mult_46_n723), .B2(mult_46_n721), .A(
        mult_46_n737), .ZN(mult_46_n736) );
  INV_X1 mult_46_U559 ( .A(mult_46_n736), .ZN(mult_46_n352) );
  XNOR2_X1 mult_46_U558 ( .A(A1[11]), .B(mult_46_n643), .ZN(mult_46_n734) );
  OAI22_X1 mult_46_U557 ( .A1(mult_46_n734), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n735), .ZN(mult_46_n353) );
  XNOR2_X1 mult_46_U556 ( .A(A1[10]), .B(mult_46_n643), .ZN(mult_46_n733) );
  OAI22_X1 mult_46_U555 ( .A1(mult_46_n733), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n734), .ZN(mult_46_n354) );
  XNOR2_X1 mult_46_U554 ( .A(A1[9]), .B(mult_46_n643), .ZN(mult_46_n732) );
  OAI22_X1 mult_46_U553 ( .A1(mult_46_n732), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n733), .ZN(mult_46_n355) );
  XNOR2_X1 mult_46_U552 ( .A(A1[8]), .B(mult_46_n643), .ZN(mult_46_n731) );
  OAI22_X1 mult_46_U551 ( .A1(mult_46_n731), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n732), .ZN(mult_46_n356) );
  XNOR2_X1 mult_46_U550 ( .A(A1[7]), .B(mult_46_n643), .ZN(mult_46_n730) );
  OAI22_X1 mult_46_U549 ( .A1(mult_46_n730), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n731), .ZN(mult_46_n357) );
  XNOR2_X1 mult_46_U548 ( .A(A1[6]), .B(mult_46_n643), .ZN(mult_46_n729) );
  OAI22_X1 mult_46_U547 ( .A1(mult_46_n729), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n730), .ZN(mult_46_n358) );
  XNOR2_X1 mult_46_U546 ( .A(A1[5]), .B(mult_46_n643), .ZN(mult_46_n728) );
  OAI22_X1 mult_46_U545 ( .A1(mult_46_n728), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n729), .ZN(mult_46_n359) );
  XNOR2_X1 mult_46_U544 ( .A(A1[4]), .B(mult_46_n643), .ZN(mult_46_n727) );
  OAI22_X1 mult_46_U543 ( .A1(mult_46_n727), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n728), .ZN(mult_46_n360) );
  XNOR2_X1 mult_46_U542 ( .A(A1[3]), .B(mult_46_n643), .ZN(mult_46_n726) );
  OAI22_X1 mult_46_U541 ( .A1(mult_46_n726), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n727), .ZN(mult_46_n361) );
  XNOR2_X1 mult_46_U540 ( .A(A1[2]), .B(mult_46_n643), .ZN(mult_46_n725) );
  OAI22_X1 mult_46_U539 ( .A1(mult_46_n725), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n726), .ZN(mult_46_n362) );
  XNOR2_X1 mult_46_U538 ( .A(A1[1]), .B(mult_46_n643), .ZN(mult_46_n724) );
  OAI22_X1 mult_46_U537 ( .A1(mult_46_n724), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n725), .ZN(mult_46_n363) );
  XNOR2_X1 mult_46_U536 ( .A(n180), .B(A1[0]), .ZN(mult_46_n722) );
  OAI22_X1 mult_46_U535 ( .A1(mult_46_n722), .A2(mult_46_n723), .B1(
        mult_46_n721), .B2(mult_46_n724), .ZN(mult_46_n364) );
  NOR2_X1 mult_46_U534 ( .A1(mult_46_n686), .A2(mult_46_n721), .ZN(
        mult_46_n365) );
  AOI21_X1 mult_46_U533 ( .B1(mult_46_n706), .B2(mult_46_n704), .A(
        mult_46_n720), .ZN(mult_46_n719) );
  INV_X1 mult_46_U532 ( .A(mult_46_n719), .ZN(mult_46_n366) );
  XNOR2_X1 mult_46_U531 ( .A(A1[11]), .B(mult_46_n641), .ZN(mult_46_n717) );
  OAI22_X1 mult_46_U530 ( .A1(mult_46_n717), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n718), .ZN(mult_46_n367) );
  XNOR2_X1 mult_46_U529 ( .A(A1[10]), .B(mult_46_n641), .ZN(mult_46_n716) );
  OAI22_X1 mult_46_U528 ( .A1(mult_46_n716), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n717), .ZN(mult_46_n368) );
  XNOR2_X1 mult_46_U527 ( .A(A1[9]), .B(mult_46_n641), .ZN(mult_46_n715) );
  OAI22_X1 mult_46_U526 ( .A1(mult_46_n715), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n716), .ZN(mult_46_n369) );
  XNOR2_X1 mult_46_U525 ( .A(A1[8]), .B(mult_46_n641), .ZN(mult_46_n714) );
  OAI22_X1 mult_46_U524 ( .A1(mult_46_n714), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n715), .ZN(mult_46_n370) );
  XNOR2_X1 mult_46_U523 ( .A(A1[7]), .B(mult_46_n641), .ZN(mult_46_n713) );
  OAI22_X1 mult_46_U522 ( .A1(mult_46_n713), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n714), .ZN(mult_46_n371) );
  XNOR2_X1 mult_46_U521 ( .A(A1[6]), .B(mult_46_n641), .ZN(mult_46_n712) );
  OAI22_X1 mult_46_U520 ( .A1(mult_46_n712), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n713), .ZN(mult_46_n372) );
  XNOR2_X1 mult_46_U519 ( .A(A1[5]), .B(mult_46_n641), .ZN(mult_46_n711) );
  OAI22_X1 mult_46_U518 ( .A1(mult_46_n711), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n712), .ZN(mult_46_n373) );
  XNOR2_X1 mult_46_U517 ( .A(A1[4]), .B(mult_46_n641), .ZN(mult_46_n710) );
  OAI22_X1 mult_46_U516 ( .A1(mult_46_n710), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n711), .ZN(mult_46_n374) );
  XNOR2_X1 mult_46_U515 ( .A(A1[3]), .B(mult_46_n641), .ZN(mult_46_n709) );
  OAI22_X1 mult_46_U514 ( .A1(mult_46_n709), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n710), .ZN(mult_46_n375) );
  XNOR2_X1 mult_46_U513 ( .A(A1[2]), .B(mult_46_n641), .ZN(mult_46_n708) );
  OAI22_X1 mult_46_U512 ( .A1(mult_46_n708), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n709), .ZN(mult_46_n376) );
  XNOR2_X1 mult_46_U511 ( .A(A1[1]), .B(mult_46_n641), .ZN(mult_46_n707) );
  OAI22_X1 mult_46_U510 ( .A1(mult_46_n707), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n708), .ZN(mult_46_n377) );
  XNOR2_X1 mult_46_U509 ( .A(mult_46_n641), .B(A1[0]), .ZN(mult_46_n705) );
  OAI22_X1 mult_46_U508 ( .A1(mult_46_n705), .A2(mult_46_n706), .B1(
        mult_46_n704), .B2(mult_46_n707), .ZN(mult_46_n378) );
  NOR2_X1 mult_46_U507 ( .A1(mult_46_n686), .A2(mult_46_n704), .ZN(
        mult_46_n379) );
  AOI21_X1 mult_46_U506 ( .B1(mult_46_n689), .B2(mult_46_n687), .A(
        mult_46_n703), .ZN(mult_46_n702) );
  INV_X1 mult_46_U505 ( .A(mult_46_n702), .ZN(mult_46_n380) );
  XNOR2_X1 mult_46_U504 ( .A(A1[11]), .B(mult_46_n639), .ZN(mult_46_n700) );
  OAI22_X1 mult_46_U503 ( .A1(mult_46_n700), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n701), .ZN(mult_46_n381) );
  OAI22_X1 mult_46_U502 ( .A1(mult_46_n699), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n700), .ZN(mult_46_n382) );
  XNOR2_X1 mult_46_U501 ( .A(A1[8]), .B(mult_46_n639), .ZN(mult_46_n697) );
  OAI22_X1 mult_46_U500 ( .A1(mult_46_n697), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n698), .ZN(mult_46_n384) );
  XNOR2_X1 mult_46_U499 ( .A(A1[7]), .B(mult_46_n639), .ZN(mult_46_n696) );
  OAI22_X1 mult_46_U498 ( .A1(mult_46_n696), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n697), .ZN(mult_46_n385) );
  XNOR2_X1 mult_46_U497 ( .A(A1[6]), .B(mult_46_n639), .ZN(mult_46_n695) );
  OAI22_X1 mult_46_U496 ( .A1(mult_46_n695), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n696), .ZN(mult_46_n386) );
  XNOR2_X1 mult_46_U495 ( .A(A1[5]), .B(mult_46_n639), .ZN(mult_46_n694) );
  OAI22_X1 mult_46_U494 ( .A1(mult_46_n694), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n695), .ZN(mult_46_n387) );
  XNOR2_X1 mult_46_U493 ( .A(A1[4]), .B(mult_46_n639), .ZN(mult_46_n693) );
  OAI22_X1 mult_46_U492 ( .A1(mult_46_n693), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n694), .ZN(mult_46_n388) );
  XNOR2_X1 mult_46_U491 ( .A(A1[3]), .B(mult_46_n639), .ZN(mult_46_n692) );
  OAI22_X1 mult_46_U490 ( .A1(mult_46_n692), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n693), .ZN(mult_46_n389) );
  XNOR2_X1 mult_46_U489 ( .A(A1[2]), .B(mult_46_n639), .ZN(mult_46_n691) );
  OAI22_X1 mult_46_U488 ( .A1(mult_46_n691), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n692), .ZN(mult_46_n390) );
  XNOR2_X1 mult_46_U487 ( .A(A1[1]), .B(mult_46_n639), .ZN(mult_46_n690) );
  OAI22_X1 mult_46_U486 ( .A1(mult_46_n690), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n691), .ZN(mult_46_n391) );
  XNOR2_X1 mult_46_U485 ( .A(n176), .B(A1[0]), .ZN(mult_46_n688) );
  OAI22_X1 mult_46_U484 ( .A1(mult_46_n688), .A2(mult_46_n689), .B1(
        mult_46_n687), .B2(mult_46_n690), .ZN(mult_46_n392) );
  NOR2_X1 mult_46_U483 ( .A1(mult_46_n686), .A2(mult_46_n687), .ZN(
        mult_46_n393) );
  AOI21_X1 mult_46_U482 ( .B1(mult_46_n670), .B2(mult_46_n671), .A(
        mult_46_n685), .ZN(mult_46_n684) );
  INV_X1 mult_46_U481 ( .A(mult_46_n684), .ZN(mult_46_n394) );
  XNOR2_X1 mult_46_U480 ( .A(A1[11]), .B(mult_46_n637), .ZN(mult_46_n682) );
  OAI22_X1 mult_46_U479 ( .A1(mult_46_n682), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n683), .ZN(mult_46_n395) );
  XNOR2_X1 mult_46_U478 ( .A(A1[10]), .B(mult_46_n637), .ZN(mult_46_n681) );
  OAI22_X1 mult_46_U477 ( .A1(mult_46_n681), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n682), .ZN(mult_46_n396) );
  XNOR2_X1 mult_46_U476 ( .A(A1[9]), .B(mult_46_n637), .ZN(mult_46_n680) );
  OAI22_X1 mult_46_U475 ( .A1(mult_46_n680), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n681), .ZN(mult_46_n397) );
  XNOR2_X1 mult_46_U474 ( .A(A1[8]), .B(mult_46_n637), .ZN(mult_46_n679) );
  OAI22_X1 mult_46_U473 ( .A1(mult_46_n679), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n680), .ZN(mult_46_n398) );
  XNOR2_X1 mult_46_U472 ( .A(A1[7]), .B(mult_46_n637), .ZN(mult_46_n678) );
  OAI22_X1 mult_46_U471 ( .A1(mult_46_n678), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n679), .ZN(mult_46_n399) );
  XNOR2_X1 mult_46_U470 ( .A(A1[6]), .B(mult_46_n637), .ZN(mult_46_n677) );
  OAI22_X1 mult_46_U469 ( .A1(mult_46_n677), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n678), .ZN(mult_46_n400) );
  XNOR2_X1 mult_46_U468 ( .A(A1[5]), .B(mult_46_n637), .ZN(mult_46_n676) );
  OAI22_X1 mult_46_U467 ( .A1(mult_46_n676), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n677), .ZN(mult_46_n401) );
  XNOR2_X1 mult_46_U466 ( .A(A1[4]), .B(mult_46_n637), .ZN(mult_46_n675) );
  OAI22_X1 mult_46_U465 ( .A1(mult_46_n675), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n676), .ZN(mult_46_n402) );
  XNOR2_X1 mult_46_U464 ( .A(A1[3]), .B(mult_46_n637), .ZN(mult_46_n674) );
  OAI22_X1 mult_46_U463 ( .A1(mult_46_n674), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n675), .ZN(mult_46_n403) );
  XNOR2_X1 mult_46_U462 ( .A(A1[2]), .B(mult_46_n637), .ZN(mult_46_n673) );
  OAI22_X1 mult_46_U461 ( .A1(mult_46_n673), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n674), .ZN(mult_46_n404) );
  XNOR2_X1 mult_46_U460 ( .A(A1[1]), .B(mult_46_n637), .ZN(mult_46_n672) );
  OAI22_X1 mult_46_U459 ( .A1(mult_46_n672), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n673), .ZN(mult_46_n405) );
  XNOR2_X1 mult_46_U458 ( .A(mult_46_n637), .B(A1[0]), .ZN(mult_46_n669) );
  OAI22_X1 mult_46_U457 ( .A1(mult_46_n669), .A2(mult_46_n670), .B1(
        mult_46_n671), .B2(mult_46_n672), .ZN(mult_46_n406) );
  XOR2_X1 mult_46_U456 ( .A(A1[13]), .B(mult_46_n636), .Z(mult_46_n667) );
  AOI21_X1 mult_46_U455 ( .B1(mult_46_n655), .B2(mult_46_n657), .A(
        mult_46_n667), .ZN(mult_46_n668) );
  INV_X1 mult_46_U454 ( .A(mult_46_n668), .ZN(mult_46_n408) );
  XNOR2_X1 mult_46_U453 ( .A(A1[12]), .B(mult_46_n635), .ZN(mult_46_n666) );
  OAI22_X1 mult_46_U452 ( .A1(mult_46_n666), .A2(mult_46_n655), .B1(
        mult_46_n667), .B2(mult_46_n657), .ZN(mult_46_n409) );
  XNOR2_X1 mult_46_U451 ( .A(A1[11]), .B(mult_46_n635), .ZN(mult_46_n665) );
  OAI22_X1 mult_46_U450 ( .A1(mult_46_n665), .A2(mult_46_n655), .B1(
        mult_46_n666), .B2(mult_46_n657), .ZN(mult_46_n410) );
  XNOR2_X1 mult_46_U449 ( .A(A1[10]), .B(mult_46_n635), .ZN(mult_46_n664) );
  OAI22_X1 mult_46_U448 ( .A1(mult_46_n664), .A2(mult_46_n655), .B1(
        mult_46_n665), .B2(mult_46_n657), .ZN(mult_46_n411) );
  XNOR2_X1 mult_46_U447 ( .A(A1[9]), .B(mult_46_n635), .ZN(mult_46_n663) );
  OAI22_X1 mult_46_U446 ( .A1(mult_46_n663), .A2(mult_46_n655), .B1(
        mult_46_n664), .B2(mult_46_n657), .ZN(mult_46_n412) );
  XNOR2_X1 mult_46_U445 ( .A(A1[8]), .B(mult_46_n635), .ZN(mult_46_n662) );
  OAI22_X1 mult_46_U444 ( .A1(mult_46_n662), .A2(mult_46_n655), .B1(
        mult_46_n663), .B2(mult_46_n657), .ZN(mult_46_n413) );
  XNOR2_X1 mult_46_U443 ( .A(A1[7]), .B(mult_46_n635), .ZN(mult_46_n661) );
  OAI22_X1 mult_46_U442 ( .A1(mult_46_n661), .A2(mult_46_n655), .B1(
        mult_46_n662), .B2(mult_46_n657), .ZN(mult_46_n414) );
  XNOR2_X1 mult_46_U441 ( .A(A1[6]), .B(mult_46_n635), .ZN(mult_46_n660) );
  OAI22_X1 mult_46_U440 ( .A1(mult_46_n660), .A2(mult_46_n655), .B1(
        mult_46_n661), .B2(mult_46_n657), .ZN(mult_46_n415) );
  XNOR2_X1 mult_46_U439 ( .A(A1[5]), .B(mult_46_n635), .ZN(mult_46_n659) );
  OAI22_X1 mult_46_U438 ( .A1(mult_46_n659), .A2(mult_46_n655), .B1(
        mult_46_n660), .B2(mult_46_n657), .ZN(mult_46_n416) );
  XNOR2_X1 mult_46_U437 ( .A(A1[4]), .B(mult_46_n635), .ZN(mult_46_n658) );
  OAI22_X1 mult_46_U436 ( .A1(mult_46_n658), .A2(mult_46_n655), .B1(
        mult_46_n659), .B2(mult_46_n657), .ZN(mult_46_n417) );
  XNOR2_X1 mult_46_U435 ( .A(A1[3]), .B(mult_46_n635), .ZN(mult_46_n656) );
  OAI22_X1 mult_46_U434 ( .A1(mult_46_n656), .A2(mult_46_n655), .B1(
        mult_46_n658), .B2(mult_46_n657), .ZN(mult_46_n418) );
  OAI22_X1 mult_46_U433 ( .A1(mult_46_n654), .A2(mult_46_n655), .B1(
        mult_46_n656), .B2(mult_46_n657), .ZN(mult_46_n419) );
  OAI21_X1 mult_46_U432 ( .B1(mult_46_n651), .B2(mult_46_n652), .A(
        mult_46_n653), .ZN(mult_46_n650) );
  XOR2_X1 mult_46_U431 ( .A(mult_46_n650), .B(mult_46_n136), .Z(mult_46_n649)
         );
  XNOR2_X1 mult_46_U430 ( .A(mult_46_n162), .B(mult_46_n649), .ZN(temp1_26_)
         );
  INV_X1 mult_46_U429 ( .A(n182), .ZN(mult_46_n646) );
  INV_X1 mult_46_U428 ( .A(n180), .ZN(mult_46_n644) );
  INV_X1 mult_46_U427 ( .A(n178), .ZN(mult_46_n642) );
  INV_X1 mult_46_U426 ( .A(n176), .ZN(mult_46_n640) );
  XOR2_X2 mult_46_U425 ( .A(reg1[12]), .B(mult_46_n646), .Z(mult_46_n755) );
  XOR2_X2 mult_46_U424 ( .A(reg1[10]), .B(mult_46_n644), .Z(mult_46_n738) );
  XOR2_X2 mult_46_U423 ( .A(reg1[8]), .B(mult_46_n642), .Z(mult_46_n721) );
  XOR2_X2 mult_46_U422 ( .A(reg1[6]), .B(mult_46_n640), .Z(mult_46_n704) );
  XOR2_X2 mult_46_U421 ( .A(reg1[4]), .B(mult_46_n638), .Z(mult_46_n687) );
  INV_X1 mult_46_U420 ( .A(reg1[0]), .ZN(mult_46_n657) );
  INV_X1 mult_46_U419 ( .A(mult_46_n805), .ZN(mult_46_n671) );
  INV_X1 mult_46_U418 ( .A(n184), .ZN(mult_46_n648) );
  INV_X1 mult_46_U417 ( .A(n172), .ZN(mult_46_n636) );
  INV_X1 mult_46_U416 ( .A(n174), .ZN(mult_46_n638) );
  INV_X1 mult_46_U415 ( .A(mult_46_n648), .ZN(mult_46_n647) );
  INV_X1 mult_46_U414 ( .A(mult_46_n646), .ZN(mult_46_n645) );
  INV_X1 mult_46_U413 ( .A(mult_46_n644), .ZN(mult_46_n643) );
  INV_X1 mult_46_U412 ( .A(mult_46_n642), .ZN(mult_46_n641) );
  INV_X1 mult_46_U411 ( .A(mult_46_n640), .ZN(mult_46_n639) );
  INV_X1 mult_46_U410 ( .A(mult_46_n636), .ZN(mult_46_n635) );
  INV_X1 mult_46_U409 ( .A(mult_46_n638), .ZN(mult_46_n637) );
  HA_X1 mult_46_U145 ( .A(mult_46_n406), .B(mult_46_n419), .CO(mult_46_n315), 
        .S(mult_46_n316) );
  FA_X1 mult_46_U144 ( .A(mult_46_n418), .B(mult_46_n393), .CI(mult_46_n405), 
        .CO(mult_46_n313), .S(mult_46_n314) );
  HA_X1 mult_46_U143 ( .A(mult_46_n321), .B(mult_46_n392), .CO(mult_46_n311), 
        .S(mult_46_n312) );
  FA_X1 mult_46_U142 ( .A(mult_46_n404), .B(mult_46_n417), .CI(mult_46_n312), 
        .CO(mult_46_n309), .S(mult_46_n310) );
  FA_X1 mult_46_U141 ( .A(mult_46_n416), .B(mult_46_n379), .CI(mult_46_n403), 
        .CO(mult_46_n307), .S(mult_46_n308) );
  FA_X1 mult_46_U140 ( .A(mult_46_n311), .B(mult_46_n391), .CI(mult_46_n308), 
        .CO(mult_46_n305), .S(mult_46_n306) );
  HA_X1 mult_46_U139 ( .A(mult_46_n320), .B(mult_46_n378), .CO(mult_46_n303), 
        .S(mult_46_n304) );
  FA_X1 mult_46_U138 ( .A(mult_46_n390), .B(mult_46_n415), .CI(mult_46_n402), 
        .CO(mult_46_n301), .S(mult_46_n302) );
  FA_X1 mult_46_U137 ( .A(mult_46_n307), .B(mult_46_n304), .CI(mult_46_n302), 
        .CO(mult_46_n299), .S(mult_46_n300) );
  FA_X1 mult_46_U136 ( .A(mult_46_n389), .B(mult_46_n365), .CI(mult_46_n414), 
        .CO(mult_46_n297), .S(mult_46_n298) );
  FA_X1 mult_46_U135 ( .A(mult_46_n377), .B(mult_46_n401), .CI(mult_46_n303), 
        .CO(mult_46_n295), .S(mult_46_n296) );
  FA_X1 mult_46_U134 ( .A(mult_46_n298), .B(mult_46_n301), .CI(mult_46_n296), 
        .CO(mult_46_n293), .S(mult_46_n294) );
  HA_X1 mult_46_U133 ( .A(mult_46_n319), .B(mult_46_n364), .CO(mult_46_n291), 
        .S(mult_46_n292) );
  FA_X1 mult_46_U132 ( .A(mult_46_n376), .B(mult_46_n388), .CI(mult_46_n400), 
        .CO(mult_46_n289), .S(mult_46_n290) );
  FA_X1 mult_46_U131 ( .A(mult_46_n292), .B(mult_46_n413), .CI(mult_46_n297), 
        .CO(mult_46_n287), .S(mult_46_n288) );
  FA_X1 mult_46_U130 ( .A(mult_46_n290), .B(mult_46_n295), .CI(mult_46_n288), 
        .CO(mult_46_n285), .S(mult_46_n286) );
  FA_X1 mult_46_U129 ( .A(mult_46_n375), .B(mult_46_n351), .CI(mult_46_n412), 
        .CO(mult_46_n283), .S(mult_46_n284) );
  FA_X1 mult_46_U128 ( .A(mult_46_n363), .B(mult_46_n399), .CI(mult_46_n387), 
        .CO(mult_46_n281), .S(mult_46_n282) );
  FA_X1 mult_46_U127 ( .A(mult_46_n289), .B(mult_46_n291), .CI(mult_46_n284), 
        .CO(mult_46_n279), .S(mult_46_n280) );
  FA_X1 mult_46_U126 ( .A(mult_46_n287), .B(mult_46_n282), .CI(mult_46_n280), 
        .CO(mult_46_n277), .S(mult_46_n278) );
  HA_X1 mult_46_U125 ( .A(mult_46_n318), .B(mult_46_n350), .CO(mult_46_n275), 
        .S(mult_46_n276) );
  FA_X1 mult_46_U124 ( .A(mult_46_n362), .B(mult_46_n386), .CI(mult_46_n411), 
        .CO(mult_46_n273), .S(mult_46_n274) );
  FA_X1 mult_46_U123 ( .A(mult_46_n374), .B(mult_46_n398), .CI(mult_46_n276), 
        .CO(mult_46_n271), .S(mult_46_n272) );
  FA_X1 mult_46_U122 ( .A(mult_46_n281), .B(mult_46_n283), .CI(mult_46_n274), 
        .CO(mult_46_n269), .S(mult_46_n270) );
  FA_X1 mult_46_U121 ( .A(mult_46_n279), .B(mult_46_n272), .CI(mult_46_n270), 
        .CO(mult_46_n267), .S(mult_46_n268) );
  FA_X1 mult_46_U120 ( .A(mult_46_n361), .B(mult_46_n337), .CI(mult_46_n410), 
        .CO(mult_46_n265), .S(mult_46_n266) );
  FA_X1 mult_46_U109 ( .A(mult_46_n349), .B(mult_46_n397), .CI(mult_46_n373), 
        .CO(mult_46_n263), .S(mult_46_n264) );
  FA_X1 mult_46_U108 ( .A(mult_46_n275), .B(mult_46_n385), .CI(mult_46_n273), 
        .CO(mult_46_n261), .S(mult_46_n262) );
  FA_X1 mult_46_U107 ( .A(mult_46_n264), .B(mult_46_n266), .CI(mult_46_n271), 
        .CO(mult_46_n259), .S(mult_46_n260) );
  FA_X1 mult_46_U106 ( .A(mult_46_n262), .B(mult_46_n269), .CI(mult_46_n260), 
        .CO(mult_46_n257), .S(mult_46_n258) );
  HA_X1 mult_46_U105 ( .A(mult_46_n317), .B(mult_46_n336), .CO(mult_46_n255), 
        .S(mult_46_n256) );
  FA_X1 mult_46_U104 ( .A(mult_46_n409), .B(mult_46_n372), .CI(mult_46_n396), 
        .CO(mult_46_n253), .S(mult_46_n254) );
  FA_X1 mult_46_U103 ( .A(mult_46_n348), .B(mult_46_n384), .CI(mult_46_n360), 
        .CO(mult_46_n251), .S(mult_46_n252) );
  FA_X1 mult_46_U102 ( .A(mult_46_n265), .B(mult_46_n256), .CI(mult_46_n263), 
        .CO(mult_46_n249), .S(mult_46_n250) );
  FA_X1 mult_46_U101 ( .A(mult_46_n254), .B(mult_46_n252), .CI(mult_46_n261), 
        .CO(mult_46_n247), .S(mult_46_n248) );
  FA_X1 mult_46_U100 ( .A(mult_46_n259), .B(mult_46_n250), .CI(mult_46_n248), 
        .CO(mult_46_n245), .S(mult_46_n246) );
  FA_X1 mult_46_U97 ( .A(mult_46_n395), .B(mult_46_n359), .CI(mult_46_n408), 
        .CO(mult_46_n241), .S(mult_46_n242) );
  FA_X1 mult_46_U96 ( .A(mult_46_n335), .B(mult_46_n371), .CI(mult_46_n255), 
        .CO(mult_46_n239), .S(mult_46_n240) );
  FA_X1 mult_46_U95 ( .A(mult_46_n253), .B(mult_46_n244), .CI(mult_46_n251), 
        .CO(mult_46_n237), .S(mult_46_n238) );
  FA_X1 mult_46_U94 ( .A(mult_46_n240), .B(mult_46_n242), .CI(mult_46_n249), 
        .CO(mult_46_n235), .S(mult_46_n236) );
  FA_X1 mult_46_U93 ( .A(mult_46_n247), .B(mult_46_n238), .CI(mult_46_n236), 
        .CO(mult_46_n233), .S(mult_46_n234) );
  FA_X1 mult_46_U91 ( .A(mult_46_n382), .B(mult_46_n346), .CI(mult_46_n232), 
        .CO(mult_46_n229), .S(mult_46_n230) );
  FA_X1 mult_46_U90 ( .A(mult_46_n334), .B(mult_46_n370), .CI(mult_46_n358), 
        .CO(mult_46_n227), .S(mult_46_n228) );
  FA_X1 mult_46_U89 ( .A(mult_46_n241), .B(mult_46_n243), .CI(mult_46_n239), 
        .CO(mult_46_n225), .S(mult_46_n226) );
  FA_X1 mult_46_U88 ( .A(mult_46_n230), .B(mult_46_n228), .CI(mult_46_n237), 
        .CO(mult_46_n223), .S(mult_46_n224) );
  FA_X1 mult_46_U87 ( .A(mult_46_n235), .B(mult_46_n226), .CI(mult_46_n224), 
        .CO(mult_46_n221), .S(mult_46_n222) );
  FA_X1 mult_46_U86 ( .A(mult_46_n231), .B(mult_46_n333), .CI(mult_46_n394), 
        .CO(mult_46_n219), .S(mult_46_n220) );
  FA_X1 mult_46_U85 ( .A(mult_46_n345), .B(mult_46_n381), .CI(mult_46_n357), 
        .CO(mult_46_n217), .S(mult_46_n218) );
  FA_X1 mult_46_U84 ( .A(mult_46_n229), .B(mult_46_n369), .CI(mult_46_n227), 
        .CO(mult_46_n215), .S(mult_46_n216) );
  FA_X1 mult_46_U83 ( .A(mult_46_n220), .B(mult_46_n218), .CI(mult_46_n225), 
        .CO(mult_46_n213), .S(mult_46_n214) );
  FA_X1 mult_46_U82 ( .A(mult_46_n223), .B(mult_46_n216), .CI(mult_46_n214), 
        .CO(mult_46_n211), .S(mult_46_n212) );
  FA_X1 mult_46_U80 ( .A(mult_46_n368), .B(mult_46_n344), .CI(mult_46_n210), 
        .CO(mult_46_n207), .S(mult_46_n208) );
  FA_X1 mult_46_U79 ( .A(mult_46_n332), .B(mult_46_n356), .CI(mult_46_n219), 
        .CO(mult_46_n205), .S(mult_46_n206) );
  FA_X1 mult_46_U78 ( .A(mult_46_n208), .B(mult_46_n217), .CI(mult_46_n215), 
        .CO(mult_46_n203), .S(mult_46_n204) );
  FA_X1 mult_46_U77 ( .A(mult_46_n213), .B(mult_46_n206), .CI(mult_46_n204), 
        .CO(mult_46_n201), .S(mult_46_n202) );
  FA_X1 mult_46_U76 ( .A(mult_46_n209), .B(mult_46_n331), .CI(mult_46_n380), 
        .CO(mult_46_n199), .S(mult_46_n200) );
  FA_X1 mult_46_U75 ( .A(mult_46_n355), .B(mult_46_n343), .CI(mult_46_n367), 
        .CO(mult_46_n197), .S(mult_46_n198) );
  FA_X1 mult_46_U74 ( .A(mult_46_n198), .B(mult_46_n207), .CI(mult_46_n200), 
        .CO(mult_46_n195), .S(mult_46_n196) );
  FA_X1 mult_46_U73 ( .A(mult_46_n203), .B(mult_46_n205), .CI(mult_46_n196), 
        .CO(mult_46_n193), .S(mult_46_n194) );
  FA_X1 mult_46_U71 ( .A(mult_46_n330), .B(mult_46_n342), .CI(mult_46_n192), 
        .CO(mult_46_n189), .S(mult_46_n190) );
  FA_X1 mult_46_U70 ( .A(mult_46_n199), .B(mult_46_n354), .CI(mult_46_n197), 
        .CO(mult_46_n187), .S(mult_46_n188) );
  FA_X1 mult_46_U69 ( .A(mult_46_n188), .B(mult_46_n190), .CI(mult_46_n195), 
        .CO(mult_46_n185), .S(mult_46_n186) );
  FA_X1 mult_46_U68 ( .A(mult_46_n191), .B(mult_46_n329), .CI(mult_46_n366), 
        .CO(mult_46_n183), .S(mult_46_n184) );
  FA_X1 mult_46_U67 ( .A(mult_46_n341), .B(mult_46_n353), .CI(mult_46_n189), 
        .CO(mult_46_n181), .S(mult_46_n182) );
  FA_X1 mult_46_U66 ( .A(mult_46_n187), .B(mult_46_n184), .CI(mult_46_n182), 
        .CO(mult_46_n179), .S(mult_46_n180) );
  FA_X1 mult_46_U64 ( .A(mult_46_n328), .B(mult_46_n340), .CI(mult_46_n178), 
        .CO(mult_46_n175), .S(mult_46_n176) );
  FA_X1 mult_46_U63 ( .A(mult_46_n176), .B(mult_46_n183), .CI(mult_46_n181), 
        .CO(mult_46_n173), .S(mult_46_n174) );
  FA_X1 mult_46_U62 ( .A(mult_46_n327), .B(mult_46_n177), .CI(mult_46_n352), 
        .CO(mult_46_n171), .S(mult_46_n172) );
  FA_X1 mult_46_U61 ( .A(mult_46_n175), .B(mult_46_n339), .CI(mult_46_n172), 
        .CO(mult_46_n169), .S(mult_46_n170) );
  FA_X1 mult_46_U59 ( .A(mult_46_n168), .B(mult_46_n326), .CI(mult_46_n171), 
        .CO(mult_46_n165), .S(mult_46_n166) );
  FA_X1 mult_46_U58 ( .A(mult_46_n325), .B(mult_46_n167), .CI(mult_46_n338), 
        .CO(mult_46_n163), .S(mult_46_n164) );
  FA_X1 mult_46_U44 ( .A(mult_46_n246), .B(mult_46_n257), .CI(mult_46_n149), 
        .CO(mult_46_n148), .S(temp1_13_) );
  FA_X1 mult_46_U43 ( .A(mult_46_n234), .B(mult_46_n245), .CI(mult_46_n148), 
        .CO(mult_46_n147), .S(temp1_14_) );
  FA_X1 mult_46_U42 ( .A(mult_46_n222), .B(mult_46_n233), .CI(mult_46_n147), 
        .CO(mult_46_n146), .S(temp1_15_) );
  FA_X1 mult_46_U41 ( .A(mult_46_n212), .B(mult_46_n221), .CI(mult_46_n146), 
        .CO(mult_46_n145), .S(temp1_16_) );
  FA_X1 mult_46_U40 ( .A(mult_46_n202), .B(mult_46_n211), .CI(mult_46_n145), 
        .CO(mult_46_n144), .S(temp1_17_) );
  FA_X1 mult_46_U39 ( .A(mult_46_n194), .B(mult_46_n201), .CI(mult_46_n144), 
        .CO(mult_46_n143), .S(temp1_18_) );
  FA_X1 mult_46_U38 ( .A(mult_46_n186), .B(mult_46_n193), .CI(mult_46_n143), 
        .CO(mult_46_n142), .S(temp1_19_) );
  FA_X1 mult_46_U37 ( .A(mult_46_n180), .B(mult_46_n185), .CI(mult_46_n142), 
        .CO(mult_46_n141), .S(temp1_20_) );
  FA_X1 mult_46_U30 ( .A(mult_46_n174), .B(mult_46_n179), .CI(mult_46_n141), 
        .CO(mult_46_n140), .S(temp1_21_) );
  FA_X1 mult_46_U20 ( .A(mult_46_n170), .B(mult_46_n173), .CI(mult_46_n140), 
        .CO(mult_46_n139), .S(temp1_22_) );
  FA_X1 mult_46_U10 ( .A(mult_46_n166), .B(mult_46_n169), .CI(mult_46_n139), 
        .CO(mult_46_n138), .S(temp1_23_) );
  FA_X1 mult_46_U9 ( .A(mult_46_n165), .B(mult_46_n164), .CI(mult_46_n138), 
        .CO(mult_46_n137), .S(temp1_24_) );
  FA_X1 mult_46_U8 ( .A(mult_46_n163), .B(mult_46_n162), .CI(mult_46_n137), 
        .CO(mult_46_n136), .S(temp1_25_) );
  XOR2_X1 mult_48_U698 ( .A(reg2[2]), .B(mult_48_n635), .Z(mult_48_n805) );
  NOR2_X1 mult_48_U697 ( .A1(mult_48_n636), .A2(A2[1]), .ZN(mult_48_n810) );
  INV_X1 mult_48_U696 ( .A(mult_48_n810), .ZN(mult_48_n812) );
  NAND2_X1 mult_48_U695 ( .A1(n158), .A2(mult_48_n657), .ZN(mult_48_n655) );
  XNOR2_X1 mult_48_U694 ( .A(A2[2]), .B(mult_48_n635), .ZN(mult_48_n654) );
  OAI22_X1 mult_48_U693 ( .A1(mult_48_n812), .A2(mult_48_n655), .B1(
        mult_48_n654), .B2(mult_48_n657), .ZN(mult_48_n811) );
  NAND2_X1 mult_48_U692 ( .A1(mult_48_n805), .A2(mult_48_n811), .ZN(
        mult_48_n808) );
  NAND2_X1 mult_48_U691 ( .A1(mult_48_n810), .A2(mult_48_n811), .ZN(
        mult_48_n809) );
  INV_X1 mult_48_U690 ( .A(A2[0]), .ZN(mult_48_n686) );
  MUX2_X1 mult_48_U689 ( .A(mult_48_n808), .B(mult_48_n809), .S(mult_48_n686), 
        .Z(mult_48_n807) );
  INV_X1 mult_48_U688 ( .A(mult_48_n807), .ZN(mult_48_n802) );
  XNOR2_X1 mult_48_U687 ( .A(mult_48_n638), .B(reg2[2]), .ZN(mult_48_n806) );
  NAND2_X1 mult_48_U686 ( .A1(mult_48_n671), .A2(mult_48_n806), .ZN(
        mult_48_n670) );
  NAND3_X1 mult_48_U685 ( .A1(mult_48_n805), .A2(mult_48_n686), .A3(
        mult_48_n637), .ZN(mult_48_n804) );
  OAI21_X1 mult_48_U684 ( .B1(mult_48_n638), .B2(mult_48_n670), .A(
        mult_48_n804), .ZN(mult_48_n803) );
  AOI222_X1 mult_48_U683 ( .A1(mult_48_n802), .A2(mult_48_n316), .B1(
        mult_48_n803), .B2(mult_48_n802), .C1(mult_48_n803), .C2(mult_48_n316), 
        .ZN(mult_48_n801) );
  INV_X1 mult_48_U682 ( .A(mult_48_n801), .ZN(mult_48_n800) );
  AOI222_X1 mult_48_U681 ( .A1(mult_48_n800), .A2(mult_48_n314), .B1(
        mult_48_n800), .B2(mult_48_n315), .C1(mult_48_n315), .C2(mult_48_n314), 
        .ZN(mult_48_n799) );
  INV_X1 mult_48_U680 ( .A(mult_48_n799), .ZN(mult_48_n798) );
  AOI222_X1 mult_48_U679 ( .A1(mult_48_n798), .A2(mult_48_n310), .B1(
        mult_48_n798), .B2(mult_48_n313), .C1(mult_48_n313), .C2(mult_48_n310), 
        .ZN(mult_48_n797) );
  INV_X1 mult_48_U678 ( .A(mult_48_n797), .ZN(mult_48_n796) );
  AOI222_X1 mult_48_U677 ( .A1(mult_48_n796), .A2(mult_48_n306), .B1(
        mult_48_n796), .B2(mult_48_n309), .C1(mult_48_n309), .C2(mult_48_n306), 
        .ZN(mult_48_n795) );
  INV_X1 mult_48_U676 ( .A(mult_48_n795), .ZN(mult_48_n794) );
  AOI222_X1 mult_48_U675 ( .A1(mult_48_n794), .A2(mult_48_n300), .B1(
        mult_48_n794), .B2(mult_48_n305), .C1(mult_48_n305), .C2(mult_48_n300), 
        .ZN(mult_48_n793) );
  INV_X1 mult_48_U674 ( .A(mult_48_n793), .ZN(mult_48_n792) );
  AOI222_X1 mult_48_U673 ( .A1(mult_48_n792), .A2(mult_48_n294), .B1(
        mult_48_n792), .B2(mult_48_n299), .C1(mult_48_n299), .C2(mult_48_n294), 
        .ZN(mult_48_n791) );
  INV_X1 mult_48_U672 ( .A(mult_48_n791), .ZN(mult_48_n790) );
  AOI222_X1 mult_48_U671 ( .A1(mult_48_n790), .A2(mult_48_n286), .B1(
        mult_48_n790), .B2(mult_48_n293), .C1(mult_48_n293), .C2(mult_48_n286), 
        .ZN(mult_48_n787) );
  INV_X1 mult_48_U670 ( .A(mult_48_n278), .ZN(mult_48_n788) );
  INV_X1 mult_48_U669 ( .A(mult_48_n285), .ZN(mult_48_n789) );
  OAI222_X1 mult_48_U668 ( .A1(mult_48_n787), .A2(mult_48_n788), .B1(
        mult_48_n787), .B2(mult_48_n789), .C1(mult_48_n789), .C2(mult_48_n788), 
        .ZN(mult_48_n786) );
  AOI222_X1 mult_48_U667 ( .A1(mult_48_n786), .A2(mult_48_n268), .B1(
        mult_48_n786), .B2(mult_48_n277), .C1(mult_48_n277), .C2(mult_48_n268), 
        .ZN(mult_48_n783) );
  INV_X1 mult_48_U666 ( .A(mult_48_n258), .ZN(mult_48_n784) );
  INV_X1 mult_48_U665 ( .A(mult_48_n267), .ZN(mult_48_n785) );
  OAI222_X1 mult_48_U664 ( .A1(mult_48_n783), .A2(mult_48_n784), .B1(
        mult_48_n783), .B2(mult_48_n785), .C1(mult_48_n785), .C2(mult_48_n784), 
        .ZN(mult_48_n149) );
  XOR2_X1 mult_48_U663 ( .A(A2[12]), .B(mult_48_n647), .Z(mult_48_n770) );
  XNOR2_X1 mult_48_U662 ( .A(mult_48_n648), .B(reg2[12]), .ZN(mult_48_n782) );
  NAND2_X1 mult_48_U661 ( .A1(mult_48_n755), .A2(mult_48_n782), .ZN(
        mult_48_n757) );
  INV_X1 mult_48_U660 ( .A(mult_48_n757), .ZN(mult_48_n651) );
  INV_X1 mult_48_U659 ( .A(mult_48_n755), .ZN(mult_48_n652) );
  XNOR2_X1 mult_48_U658 ( .A(A2[13]), .B(mult_48_n648), .ZN(mult_48_n653) );
  AOI22_X1 mult_48_U657 ( .A1(mult_48_n770), .A2(mult_48_n651), .B1(
        mult_48_n652), .B2(mult_48_n653), .ZN(mult_48_n162) );
  XNOR2_X1 mult_48_U656 ( .A(A2[12]), .B(mult_48_n645), .ZN(mult_48_n752) );
  XNOR2_X1 mult_48_U655 ( .A(mult_48_n646), .B(reg2[10]), .ZN(mult_48_n781) );
  NAND2_X1 mult_48_U654 ( .A1(mult_48_n738), .A2(mult_48_n781), .ZN(
        mult_48_n740) );
  XNOR2_X1 mult_48_U653 ( .A(A2[13]), .B(mult_48_n645), .ZN(mult_48_n754) );
  OAI22_X1 mult_48_U652 ( .A1(mult_48_n752), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n754), .ZN(mult_48_n167) );
  INV_X1 mult_48_U651 ( .A(mult_48_n167), .ZN(mult_48_n168) );
  XNOR2_X1 mult_48_U650 ( .A(A2[12]), .B(mult_48_n643), .ZN(mult_48_n735) );
  XNOR2_X1 mult_48_U649 ( .A(mult_48_n644), .B(reg2[8]), .ZN(mult_48_n780) );
  NAND2_X1 mult_48_U648 ( .A1(mult_48_n721), .A2(mult_48_n780), .ZN(
        mult_48_n723) );
  XNOR2_X1 mult_48_U647 ( .A(A2[13]), .B(mult_48_n643), .ZN(mult_48_n737) );
  OAI22_X1 mult_48_U646 ( .A1(mult_48_n735), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n737), .ZN(mult_48_n177) );
  INV_X1 mult_48_U645 ( .A(mult_48_n177), .ZN(mult_48_n178) );
  XNOR2_X1 mult_48_U644 ( .A(A2[12]), .B(mult_48_n641), .ZN(mult_48_n718) );
  XNOR2_X1 mult_48_U643 ( .A(mult_48_n642), .B(reg2[6]), .ZN(mult_48_n779) );
  NAND2_X1 mult_48_U642 ( .A1(mult_48_n704), .A2(mult_48_n779), .ZN(
        mult_48_n706) );
  XNOR2_X1 mult_48_U641 ( .A(A2[13]), .B(mult_48_n641), .ZN(mult_48_n720) );
  OAI22_X1 mult_48_U640 ( .A1(mult_48_n718), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n720), .ZN(mult_48_n191) );
  INV_X1 mult_48_U639 ( .A(mult_48_n191), .ZN(mult_48_n192) );
  XNOR2_X1 mult_48_U638 ( .A(A2[12]), .B(mult_48_n639), .ZN(mult_48_n701) );
  XNOR2_X1 mult_48_U637 ( .A(mult_48_n640), .B(reg2[4]), .ZN(mult_48_n778) );
  NAND2_X1 mult_48_U636 ( .A1(mult_48_n687), .A2(mult_48_n778), .ZN(
        mult_48_n689) );
  XNOR2_X1 mult_48_U635 ( .A(A2[13]), .B(mult_48_n639), .ZN(mult_48_n703) );
  OAI22_X1 mult_48_U634 ( .A1(mult_48_n701), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n703), .ZN(mult_48_n209) );
  INV_X1 mult_48_U633 ( .A(mult_48_n209), .ZN(mult_48_n210) );
  XNOR2_X1 mult_48_U632 ( .A(A2[12]), .B(mult_48_n637), .ZN(mult_48_n683) );
  XNOR2_X1 mult_48_U631 ( .A(A2[13]), .B(mult_48_n637), .ZN(mult_48_n685) );
  OAI22_X1 mult_48_U630 ( .A1(mult_48_n683), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n685), .ZN(mult_48_n231) );
  INV_X1 mult_48_U629 ( .A(mult_48_n231), .ZN(mult_48_n232) );
  XNOR2_X1 mult_48_U628 ( .A(A2[3]), .B(mult_48_n645), .ZN(mult_48_n743) );
  XNOR2_X1 mult_48_U627 ( .A(A2[4]), .B(mult_48_n645), .ZN(mult_48_n744) );
  OAI22_X1 mult_48_U626 ( .A1(mult_48_n743), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n744), .ZN(mult_48_n776) );
  XNOR2_X1 mult_48_U625 ( .A(A2[9]), .B(mult_48_n639), .ZN(mult_48_n698) );
  XNOR2_X1 mult_48_U624 ( .A(A2[10]), .B(mult_48_n639), .ZN(mult_48_n699) );
  OAI22_X1 mult_48_U623 ( .A1(mult_48_n698), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n699), .ZN(mult_48_n777) );
  OR2_X1 mult_48_U622 ( .A1(mult_48_n776), .A2(mult_48_n777), .ZN(mult_48_n243) );
  XNOR2_X1 mult_48_U621 ( .A(mult_48_n776), .B(mult_48_n777), .ZN(mult_48_n244) );
  NAND3_X1 mult_48_U620 ( .A1(mult_48_n652), .A2(mult_48_n686), .A3(n170), 
        .ZN(mult_48_n775) );
  OAI21_X1 mult_48_U619 ( .B1(mult_48_n648), .B2(mult_48_n757), .A(
        mult_48_n775), .ZN(mult_48_n317) );
  OR3_X1 mult_48_U618 ( .A1(mult_48_n738), .A2(A2[0]), .A3(mult_48_n646), .ZN(
        mult_48_n774) );
  OAI21_X1 mult_48_U617 ( .B1(mult_48_n646), .B2(mult_48_n740), .A(
        mult_48_n774), .ZN(mult_48_n318) );
  OR3_X1 mult_48_U616 ( .A1(mult_48_n721), .A2(A2[0]), .A3(mult_48_n644), .ZN(
        mult_48_n773) );
  OAI21_X1 mult_48_U615 ( .B1(mult_48_n644), .B2(mult_48_n723), .A(
        mult_48_n773), .ZN(mult_48_n319) );
  OR3_X1 mult_48_U614 ( .A1(mult_48_n704), .A2(A2[0]), .A3(mult_48_n642), .ZN(
        mult_48_n772) );
  OAI21_X1 mult_48_U613 ( .B1(mult_48_n642), .B2(mult_48_n706), .A(
        mult_48_n772), .ZN(mult_48_n320) );
  OR3_X1 mult_48_U612 ( .A1(mult_48_n687), .A2(A2[0]), .A3(mult_48_n640), .ZN(
        mult_48_n771) );
  OAI21_X1 mult_48_U611 ( .B1(mult_48_n640), .B2(mult_48_n689), .A(
        mult_48_n771), .ZN(mult_48_n321) );
  XNOR2_X1 mult_48_U610 ( .A(A2[11]), .B(mult_48_n647), .ZN(mult_48_n768) );
  INV_X1 mult_48_U609 ( .A(mult_48_n770), .ZN(mult_48_n769) );
  OAI22_X1 mult_48_U608 ( .A1(mult_48_n768), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n769), .ZN(mult_48_n325) );
  XNOR2_X1 mult_48_U607 ( .A(A2[10]), .B(mult_48_n647), .ZN(mult_48_n767) );
  OAI22_X1 mult_48_U606 ( .A1(mult_48_n767), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n768), .ZN(mult_48_n326) );
  XNOR2_X1 mult_48_U605 ( .A(A2[9]), .B(mult_48_n647), .ZN(mult_48_n766) );
  OAI22_X1 mult_48_U604 ( .A1(mult_48_n766), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n767), .ZN(mult_48_n327) );
  XNOR2_X1 mult_48_U603 ( .A(A2[8]), .B(mult_48_n647), .ZN(mult_48_n765) );
  OAI22_X1 mult_48_U602 ( .A1(mult_48_n765), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n766), .ZN(mult_48_n328) );
  XNOR2_X1 mult_48_U601 ( .A(A2[7]), .B(mult_48_n647), .ZN(mult_48_n764) );
  OAI22_X1 mult_48_U600 ( .A1(mult_48_n764), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n765), .ZN(mult_48_n329) );
  XNOR2_X1 mult_48_U599 ( .A(A2[6]), .B(mult_48_n647), .ZN(mult_48_n763) );
  OAI22_X1 mult_48_U598 ( .A1(mult_48_n763), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n764), .ZN(mult_48_n330) );
  XNOR2_X1 mult_48_U597 ( .A(A2[5]), .B(mult_48_n647), .ZN(mult_48_n762) );
  OAI22_X1 mult_48_U596 ( .A1(mult_48_n762), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n763), .ZN(mult_48_n331) );
  XNOR2_X1 mult_48_U595 ( .A(A2[4]), .B(mult_48_n647), .ZN(mult_48_n761) );
  OAI22_X1 mult_48_U594 ( .A1(mult_48_n761), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n762), .ZN(mult_48_n332) );
  XNOR2_X1 mult_48_U593 ( .A(A2[3]), .B(mult_48_n647), .ZN(mult_48_n760) );
  OAI22_X1 mult_48_U592 ( .A1(mult_48_n760), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n761), .ZN(mult_48_n333) );
  XNOR2_X1 mult_48_U591 ( .A(A2[2]), .B(mult_48_n647), .ZN(mult_48_n759) );
  OAI22_X1 mult_48_U590 ( .A1(mult_48_n759), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n760), .ZN(mult_48_n334) );
  XNOR2_X1 mult_48_U589 ( .A(A2[1]), .B(mult_48_n647), .ZN(mult_48_n758) );
  OAI22_X1 mult_48_U588 ( .A1(mult_48_n758), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n759), .ZN(mult_48_n335) );
  XNOR2_X1 mult_48_U587 ( .A(n170), .B(A2[0]), .ZN(mult_48_n756) );
  OAI22_X1 mult_48_U586 ( .A1(mult_48_n756), .A2(mult_48_n757), .B1(
        mult_48_n755), .B2(mult_48_n758), .ZN(mult_48_n336) );
  NOR2_X1 mult_48_U585 ( .A1(mult_48_n686), .A2(mult_48_n755), .ZN(
        mult_48_n337) );
  AOI21_X1 mult_48_U584 ( .B1(mult_48_n740), .B2(mult_48_n738), .A(
        mult_48_n754), .ZN(mult_48_n753) );
  INV_X1 mult_48_U583 ( .A(mult_48_n753), .ZN(mult_48_n338) );
  XNOR2_X1 mult_48_U582 ( .A(A2[11]), .B(mult_48_n645), .ZN(mult_48_n751) );
  OAI22_X1 mult_48_U581 ( .A1(mult_48_n751), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n752), .ZN(mult_48_n339) );
  XNOR2_X1 mult_48_U580 ( .A(A2[10]), .B(mult_48_n645), .ZN(mult_48_n750) );
  OAI22_X1 mult_48_U579 ( .A1(mult_48_n750), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n751), .ZN(mult_48_n340) );
  XNOR2_X1 mult_48_U578 ( .A(A2[9]), .B(mult_48_n645), .ZN(mult_48_n749) );
  OAI22_X1 mult_48_U577 ( .A1(mult_48_n749), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n750), .ZN(mult_48_n341) );
  XNOR2_X1 mult_48_U576 ( .A(A2[8]), .B(mult_48_n645), .ZN(mult_48_n748) );
  OAI22_X1 mult_48_U575 ( .A1(mult_48_n748), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n749), .ZN(mult_48_n342) );
  XNOR2_X1 mult_48_U574 ( .A(A2[7]), .B(mult_48_n645), .ZN(mult_48_n747) );
  OAI22_X1 mult_48_U573 ( .A1(mult_48_n747), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n748), .ZN(mult_48_n343) );
  XNOR2_X1 mult_48_U572 ( .A(A2[6]), .B(mult_48_n645), .ZN(mult_48_n746) );
  OAI22_X1 mult_48_U571 ( .A1(mult_48_n746), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n747), .ZN(mult_48_n344) );
  XNOR2_X1 mult_48_U570 ( .A(A2[5]), .B(mult_48_n645), .ZN(mult_48_n745) );
  OAI22_X1 mult_48_U569 ( .A1(mult_48_n745), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n746), .ZN(mult_48_n345) );
  OAI22_X1 mult_48_U568 ( .A1(mult_48_n744), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n745), .ZN(mult_48_n346) );
  XNOR2_X1 mult_48_U567 ( .A(A2[2]), .B(mult_48_n645), .ZN(mult_48_n742) );
  OAI22_X1 mult_48_U566 ( .A1(mult_48_n742), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n743), .ZN(mult_48_n348) );
  XNOR2_X1 mult_48_U565 ( .A(A2[1]), .B(mult_48_n645), .ZN(mult_48_n741) );
  OAI22_X1 mult_48_U564 ( .A1(mult_48_n741), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n742), .ZN(mult_48_n349) );
  XNOR2_X1 mult_48_U563 ( .A(n168), .B(A2[0]), .ZN(mult_48_n739) );
  OAI22_X1 mult_48_U562 ( .A1(mult_48_n739), .A2(mult_48_n740), .B1(
        mult_48_n738), .B2(mult_48_n741), .ZN(mult_48_n350) );
  NOR2_X1 mult_48_U561 ( .A1(mult_48_n686), .A2(mult_48_n738), .ZN(
        mult_48_n351) );
  AOI21_X1 mult_48_U560 ( .B1(mult_48_n723), .B2(mult_48_n721), .A(
        mult_48_n737), .ZN(mult_48_n736) );
  INV_X1 mult_48_U559 ( .A(mult_48_n736), .ZN(mult_48_n352) );
  XNOR2_X1 mult_48_U558 ( .A(A2[11]), .B(mult_48_n643), .ZN(mult_48_n734) );
  OAI22_X1 mult_48_U557 ( .A1(mult_48_n734), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n735), .ZN(mult_48_n353) );
  XNOR2_X1 mult_48_U556 ( .A(A2[10]), .B(mult_48_n643), .ZN(mult_48_n733) );
  OAI22_X1 mult_48_U555 ( .A1(mult_48_n733), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n734), .ZN(mult_48_n354) );
  XNOR2_X1 mult_48_U554 ( .A(A2[9]), .B(mult_48_n643), .ZN(mult_48_n732) );
  OAI22_X1 mult_48_U553 ( .A1(mult_48_n732), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n733), .ZN(mult_48_n355) );
  XNOR2_X1 mult_48_U552 ( .A(A2[8]), .B(mult_48_n643), .ZN(mult_48_n731) );
  OAI22_X1 mult_48_U551 ( .A1(mult_48_n731), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n732), .ZN(mult_48_n356) );
  XNOR2_X1 mult_48_U550 ( .A(A2[7]), .B(mult_48_n643), .ZN(mult_48_n730) );
  OAI22_X1 mult_48_U549 ( .A1(mult_48_n730), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n731), .ZN(mult_48_n357) );
  XNOR2_X1 mult_48_U548 ( .A(A2[6]), .B(mult_48_n643), .ZN(mult_48_n729) );
  OAI22_X1 mult_48_U547 ( .A1(mult_48_n729), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n730), .ZN(mult_48_n358) );
  XNOR2_X1 mult_48_U546 ( .A(A2[5]), .B(mult_48_n643), .ZN(mult_48_n728) );
  OAI22_X1 mult_48_U545 ( .A1(mult_48_n728), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n729), .ZN(mult_48_n359) );
  XNOR2_X1 mult_48_U544 ( .A(A2[4]), .B(mult_48_n643), .ZN(mult_48_n727) );
  OAI22_X1 mult_48_U543 ( .A1(mult_48_n727), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n728), .ZN(mult_48_n360) );
  XNOR2_X1 mult_48_U542 ( .A(A2[3]), .B(mult_48_n643), .ZN(mult_48_n726) );
  OAI22_X1 mult_48_U541 ( .A1(mult_48_n726), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n727), .ZN(mult_48_n361) );
  XNOR2_X1 mult_48_U540 ( .A(A2[2]), .B(mult_48_n643), .ZN(mult_48_n725) );
  OAI22_X1 mult_48_U539 ( .A1(mult_48_n725), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n726), .ZN(mult_48_n362) );
  XNOR2_X1 mult_48_U538 ( .A(A2[1]), .B(mult_48_n643), .ZN(mult_48_n724) );
  OAI22_X1 mult_48_U537 ( .A1(mult_48_n724), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n725), .ZN(mult_48_n363) );
  XNOR2_X1 mult_48_U536 ( .A(n166), .B(A2[0]), .ZN(mult_48_n722) );
  OAI22_X1 mult_48_U535 ( .A1(mult_48_n722), .A2(mult_48_n723), .B1(
        mult_48_n721), .B2(mult_48_n724), .ZN(mult_48_n364) );
  NOR2_X1 mult_48_U534 ( .A1(mult_48_n686), .A2(mult_48_n721), .ZN(
        mult_48_n365) );
  AOI21_X1 mult_48_U533 ( .B1(mult_48_n706), .B2(mult_48_n704), .A(
        mult_48_n720), .ZN(mult_48_n719) );
  INV_X1 mult_48_U532 ( .A(mult_48_n719), .ZN(mult_48_n366) );
  XNOR2_X1 mult_48_U531 ( .A(A2[11]), .B(mult_48_n641), .ZN(mult_48_n717) );
  OAI22_X1 mult_48_U530 ( .A1(mult_48_n717), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n718), .ZN(mult_48_n367) );
  XNOR2_X1 mult_48_U529 ( .A(A2[10]), .B(mult_48_n641), .ZN(mult_48_n716) );
  OAI22_X1 mult_48_U528 ( .A1(mult_48_n716), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n717), .ZN(mult_48_n368) );
  XNOR2_X1 mult_48_U527 ( .A(A2[9]), .B(mult_48_n641), .ZN(mult_48_n715) );
  OAI22_X1 mult_48_U526 ( .A1(mult_48_n715), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n716), .ZN(mult_48_n369) );
  XNOR2_X1 mult_48_U525 ( .A(A2[8]), .B(mult_48_n641), .ZN(mult_48_n714) );
  OAI22_X1 mult_48_U524 ( .A1(mult_48_n714), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n715), .ZN(mult_48_n370) );
  XNOR2_X1 mult_48_U523 ( .A(A2[7]), .B(mult_48_n641), .ZN(mult_48_n713) );
  OAI22_X1 mult_48_U522 ( .A1(mult_48_n713), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n714), .ZN(mult_48_n371) );
  XNOR2_X1 mult_48_U521 ( .A(A2[6]), .B(mult_48_n641), .ZN(mult_48_n712) );
  OAI22_X1 mult_48_U520 ( .A1(mult_48_n712), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n713), .ZN(mult_48_n372) );
  XNOR2_X1 mult_48_U519 ( .A(A2[5]), .B(mult_48_n641), .ZN(mult_48_n711) );
  OAI22_X1 mult_48_U518 ( .A1(mult_48_n711), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n712), .ZN(mult_48_n373) );
  XNOR2_X1 mult_48_U517 ( .A(A2[4]), .B(mult_48_n641), .ZN(mult_48_n710) );
  OAI22_X1 mult_48_U516 ( .A1(mult_48_n710), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n711), .ZN(mult_48_n374) );
  XNOR2_X1 mult_48_U515 ( .A(A2[3]), .B(mult_48_n641), .ZN(mult_48_n709) );
  OAI22_X1 mult_48_U514 ( .A1(mult_48_n709), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n710), .ZN(mult_48_n375) );
  XNOR2_X1 mult_48_U513 ( .A(A2[2]), .B(mult_48_n641), .ZN(mult_48_n708) );
  OAI22_X1 mult_48_U512 ( .A1(mult_48_n708), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n709), .ZN(mult_48_n376) );
  XNOR2_X1 mult_48_U511 ( .A(A2[1]), .B(mult_48_n641), .ZN(mult_48_n707) );
  OAI22_X1 mult_48_U510 ( .A1(mult_48_n707), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n708), .ZN(mult_48_n377) );
  XNOR2_X1 mult_48_U509 ( .A(mult_48_n641), .B(A2[0]), .ZN(mult_48_n705) );
  OAI22_X1 mult_48_U508 ( .A1(mult_48_n705), .A2(mult_48_n706), .B1(
        mult_48_n704), .B2(mult_48_n707), .ZN(mult_48_n378) );
  NOR2_X1 mult_48_U507 ( .A1(mult_48_n686), .A2(mult_48_n704), .ZN(
        mult_48_n379) );
  AOI21_X1 mult_48_U506 ( .B1(mult_48_n689), .B2(mult_48_n687), .A(
        mult_48_n703), .ZN(mult_48_n702) );
  INV_X1 mult_48_U505 ( .A(mult_48_n702), .ZN(mult_48_n380) );
  XNOR2_X1 mult_48_U504 ( .A(A2[11]), .B(mult_48_n639), .ZN(mult_48_n700) );
  OAI22_X1 mult_48_U503 ( .A1(mult_48_n700), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n701), .ZN(mult_48_n381) );
  OAI22_X1 mult_48_U502 ( .A1(mult_48_n699), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n700), .ZN(mult_48_n382) );
  XNOR2_X1 mult_48_U501 ( .A(A2[8]), .B(mult_48_n639), .ZN(mult_48_n697) );
  OAI22_X1 mult_48_U500 ( .A1(mult_48_n697), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n698), .ZN(mult_48_n384) );
  XNOR2_X1 mult_48_U499 ( .A(A2[7]), .B(mult_48_n639), .ZN(mult_48_n696) );
  OAI22_X1 mult_48_U498 ( .A1(mult_48_n696), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n697), .ZN(mult_48_n385) );
  XNOR2_X1 mult_48_U497 ( .A(A2[6]), .B(mult_48_n639), .ZN(mult_48_n695) );
  OAI22_X1 mult_48_U496 ( .A1(mult_48_n695), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n696), .ZN(mult_48_n386) );
  XNOR2_X1 mult_48_U495 ( .A(A2[5]), .B(mult_48_n639), .ZN(mult_48_n694) );
  OAI22_X1 mult_48_U494 ( .A1(mult_48_n694), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n695), .ZN(mult_48_n387) );
  XNOR2_X1 mult_48_U493 ( .A(A2[4]), .B(mult_48_n639), .ZN(mult_48_n693) );
  OAI22_X1 mult_48_U492 ( .A1(mult_48_n693), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n694), .ZN(mult_48_n388) );
  XNOR2_X1 mult_48_U491 ( .A(A2[3]), .B(mult_48_n639), .ZN(mult_48_n692) );
  OAI22_X1 mult_48_U490 ( .A1(mult_48_n692), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n693), .ZN(mult_48_n389) );
  XNOR2_X1 mult_48_U489 ( .A(A2[2]), .B(mult_48_n639), .ZN(mult_48_n691) );
  OAI22_X1 mult_48_U488 ( .A1(mult_48_n691), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n692), .ZN(mult_48_n390) );
  XNOR2_X1 mult_48_U487 ( .A(A2[1]), .B(mult_48_n639), .ZN(mult_48_n690) );
  OAI22_X1 mult_48_U486 ( .A1(mult_48_n690), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n691), .ZN(mult_48_n391) );
  XNOR2_X1 mult_48_U485 ( .A(n162), .B(A2[0]), .ZN(mult_48_n688) );
  OAI22_X1 mult_48_U484 ( .A1(mult_48_n688), .A2(mult_48_n689), .B1(
        mult_48_n687), .B2(mult_48_n690), .ZN(mult_48_n392) );
  NOR2_X1 mult_48_U483 ( .A1(mult_48_n686), .A2(mult_48_n687), .ZN(
        mult_48_n393) );
  AOI21_X1 mult_48_U482 ( .B1(mult_48_n670), .B2(mult_48_n671), .A(
        mult_48_n685), .ZN(mult_48_n684) );
  INV_X1 mult_48_U481 ( .A(mult_48_n684), .ZN(mult_48_n394) );
  XNOR2_X1 mult_48_U480 ( .A(A2[11]), .B(mult_48_n637), .ZN(mult_48_n682) );
  OAI22_X1 mult_48_U479 ( .A1(mult_48_n682), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n683), .ZN(mult_48_n395) );
  XNOR2_X1 mult_48_U478 ( .A(A2[10]), .B(mult_48_n637), .ZN(mult_48_n681) );
  OAI22_X1 mult_48_U477 ( .A1(mult_48_n681), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n682), .ZN(mult_48_n396) );
  XNOR2_X1 mult_48_U476 ( .A(A2[9]), .B(mult_48_n637), .ZN(mult_48_n680) );
  OAI22_X1 mult_48_U475 ( .A1(mult_48_n680), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n681), .ZN(mult_48_n397) );
  XNOR2_X1 mult_48_U474 ( .A(A2[8]), .B(mult_48_n637), .ZN(mult_48_n679) );
  OAI22_X1 mult_48_U473 ( .A1(mult_48_n679), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n680), .ZN(mult_48_n398) );
  XNOR2_X1 mult_48_U472 ( .A(A2[7]), .B(mult_48_n637), .ZN(mult_48_n678) );
  OAI22_X1 mult_48_U471 ( .A1(mult_48_n678), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n679), .ZN(mult_48_n399) );
  XNOR2_X1 mult_48_U470 ( .A(A2[6]), .B(mult_48_n637), .ZN(mult_48_n677) );
  OAI22_X1 mult_48_U469 ( .A1(mult_48_n677), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n678), .ZN(mult_48_n400) );
  XNOR2_X1 mult_48_U468 ( .A(A2[5]), .B(mult_48_n637), .ZN(mult_48_n676) );
  OAI22_X1 mult_48_U467 ( .A1(mult_48_n676), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n677), .ZN(mult_48_n401) );
  XNOR2_X1 mult_48_U466 ( .A(A2[4]), .B(mult_48_n637), .ZN(mult_48_n675) );
  OAI22_X1 mult_48_U465 ( .A1(mult_48_n675), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n676), .ZN(mult_48_n402) );
  XNOR2_X1 mult_48_U464 ( .A(A2[3]), .B(mult_48_n637), .ZN(mult_48_n674) );
  OAI22_X1 mult_48_U463 ( .A1(mult_48_n674), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n675), .ZN(mult_48_n403) );
  XNOR2_X1 mult_48_U462 ( .A(A2[2]), .B(mult_48_n637), .ZN(mult_48_n673) );
  OAI22_X1 mult_48_U461 ( .A1(mult_48_n673), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n674), .ZN(mult_48_n404) );
  XNOR2_X1 mult_48_U460 ( .A(A2[1]), .B(mult_48_n637), .ZN(mult_48_n672) );
  OAI22_X1 mult_48_U459 ( .A1(mult_48_n672), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n673), .ZN(mult_48_n405) );
  XNOR2_X1 mult_48_U458 ( .A(mult_48_n637), .B(A2[0]), .ZN(mult_48_n669) );
  OAI22_X1 mult_48_U457 ( .A1(mult_48_n669), .A2(mult_48_n670), .B1(
        mult_48_n671), .B2(mult_48_n672), .ZN(mult_48_n406) );
  XOR2_X1 mult_48_U456 ( .A(A2[13]), .B(mult_48_n636), .Z(mult_48_n667) );
  AOI21_X1 mult_48_U455 ( .B1(mult_48_n655), .B2(mult_48_n657), .A(
        mult_48_n667), .ZN(mult_48_n668) );
  INV_X1 mult_48_U454 ( .A(mult_48_n668), .ZN(mult_48_n408) );
  XNOR2_X1 mult_48_U453 ( .A(A2[12]), .B(mult_48_n635), .ZN(mult_48_n666) );
  OAI22_X1 mult_48_U452 ( .A1(mult_48_n666), .A2(mult_48_n655), .B1(
        mult_48_n667), .B2(mult_48_n657), .ZN(mult_48_n409) );
  XNOR2_X1 mult_48_U451 ( .A(A2[11]), .B(mult_48_n635), .ZN(mult_48_n665) );
  OAI22_X1 mult_48_U450 ( .A1(mult_48_n665), .A2(mult_48_n655), .B1(
        mult_48_n666), .B2(mult_48_n657), .ZN(mult_48_n410) );
  XNOR2_X1 mult_48_U449 ( .A(A2[10]), .B(mult_48_n635), .ZN(mult_48_n664) );
  OAI22_X1 mult_48_U448 ( .A1(mult_48_n664), .A2(mult_48_n655), .B1(
        mult_48_n665), .B2(mult_48_n657), .ZN(mult_48_n411) );
  XNOR2_X1 mult_48_U447 ( .A(A2[9]), .B(mult_48_n635), .ZN(mult_48_n663) );
  OAI22_X1 mult_48_U446 ( .A1(mult_48_n663), .A2(mult_48_n655), .B1(
        mult_48_n664), .B2(mult_48_n657), .ZN(mult_48_n412) );
  XNOR2_X1 mult_48_U445 ( .A(A2[8]), .B(mult_48_n635), .ZN(mult_48_n662) );
  OAI22_X1 mult_48_U444 ( .A1(mult_48_n662), .A2(mult_48_n655), .B1(
        mult_48_n663), .B2(mult_48_n657), .ZN(mult_48_n413) );
  XNOR2_X1 mult_48_U443 ( .A(A2[7]), .B(mult_48_n635), .ZN(mult_48_n661) );
  OAI22_X1 mult_48_U442 ( .A1(mult_48_n661), .A2(mult_48_n655), .B1(
        mult_48_n662), .B2(mult_48_n657), .ZN(mult_48_n414) );
  XNOR2_X1 mult_48_U441 ( .A(A2[6]), .B(mult_48_n635), .ZN(mult_48_n660) );
  OAI22_X1 mult_48_U440 ( .A1(mult_48_n660), .A2(mult_48_n655), .B1(
        mult_48_n661), .B2(mult_48_n657), .ZN(mult_48_n415) );
  XNOR2_X1 mult_48_U439 ( .A(A2[5]), .B(mult_48_n635), .ZN(mult_48_n659) );
  OAI22_X1 mult_48_U438 ( .A1(mult_48_n659), .A2(mult_48_n655), .B1(
        mult_48_n660), .B2(mult_48_n657), .ZN(mult_48_n416) );
  XNOR2_X1 mult_48_U437 ( .A(A2[4]), .B(mult_48_n635), .ZN(mult_48_n658) );
  OAI22_X1 mult_48_U436 ( .A1(mult_48_n658), .A2(mult_48_n655), .B1(
        mult_48_n659), .B2(mult_48_n657), .ZN(mult_48_n417) );
  XNOR2_X1 mult_48_U435 ( .A(A2[3]), .B(mult_48_n635), .ZN(mult_48_n656) );
  OAI22_X1 mult_48_U434 ( .A1(mult_48_n656), .A2(mult_48_n655), .B1(
        mult_48_n658), .B2(mult_48_n657), .ZN(mult_48_n418) );
  OAI22_X1 mult_48_U433 ( .A1(mult_48_n654), .A2(mult_48_n655), .B1(
        mult_48_n656), .B2(mult_48_n657), .ZN(mult_48_n419) );
  OAI21_X1 mult_48_U432 ( .B1(mult_48_n651), .B2(mult_48_n652), .A(
        mult_48_n653), .ZN(mult_48_n650) );
  XOR2_X1 mult_48_U431 ( .A(mult_48_n650), .B(mult_48_n136), .Z(mult_48_n649)
         );
  XNOR2_X1 mult_48_U430 ( .A(mult_48_n162), .B(mult_48_n649), .ZN(temp2_26_)
         );
  INV_X1 mult_48_U429 ( .A(n168), .ZN(mult_48_n646) );
  INV_X1 mult_48_U428 ( .A(n166), .ZN(mult_48_n644) );
  INV_X1 mult_48_U427 ( .A(n164), .ZN(mult_48_n642) );
  INV_X1 mult_48_U426 ( .A(n162), .ZN(mult_48_n640) );
  XOR2_X2 mult_48_U425 ( .A(reg2[12]), .B(mult_48_n646), .Z(mult_48_n755) );
  XOR2_X2 mult_48_U424 ( .A(reg2[10]), .B(mult_48_n644), .Z(mult_48_n738) );
  XOR2_X2 mult_48_U423 ( .A(reg2[8]), .B(mult_48_n642), .Z(mult_48_n721) );
  XOR2_X2 mult_48_U422 ( .A(reg2[6]), .B(mult_48_n640), .Z(mult_48_n704) );
  XOR2_X2 mult_48_U421 ( .A(reg2[4]), .B(mult_48_n638), .Z(mult_48_n687) );
  INV_X1 mult_48_U420 ( .A(reg2[0]), .ZN(mult_48_n657) );
  INV_X1 mult_48_U419 ( .A(mult_48_n805), .ZN(mult_48_n671) );
  INV_X1 mult_48_U418 ( .A(n170), .ZN(mult_48_n648) );
  INV_X1 mult_48_U417 ( .A(n158), .ZN(mult_48_n636) );
  INV_X1 mult_48_U416 ( .A(n160), .ZN(mult_48_n638) );
  INV_X1 mult_48_U415 ( .A(mult_48_n648), .ZN(mult_48_n647) );
  INV_X1 mult_48_U414 ( .A(mult_48_n646), .ZN(mult_48_n645) );
  INV_X1 mult_48_U413 ( .A(mult_48_n644), .ZN(mult_48_n643) );
  INV_X1 mult_48_U412 ( .A(mult_48_n642), .ZN(mult_48_n641) );
  INV_X1 mult_48_U411 ( .A(mult_48_n640), .ZN(mult_48_n639) );
  INV_X1 mult_48_U410 ( .A(mult_48_n638), .ZN(mult_48_n637) );
  INV_X1 mult_48_U409 ( .A(mult_48_n636), .ZN(mult_48_n635) );
  HA_X1 mult_48_U145 ( .A(mult_48_n406), .B(mult_48_n419), .CO(mult_48_n315), 
        .S(mult_48_n316) );
  FA_X1 mult_48_U144 ( .A(mult_48_n418), .B(mult_48_n393), .CI(mult_48_n405), 
        .CO(mult_48_n313), .S(mult_48_n314) );
  HA_X1 mult_48_U143 ( .A(mult_48_n321), .B(mult_48_n392), .CO(mult_48_n311), 
        .S(mult_48_n312) );
  FA_X1 mult_48_U142 ( .A(mult_48_n404), .B(mult_48_n417), .CI(mult_48_n312), 
        .CO(mult_48_n309), .S(mult_48_n310) );
  FA_X1 mult_48_U141 ( .A(mult_48_n416), .B(mult_48_n379), .CI(mult_48_n403), 
        .CO(mult_48_n307), .S(mult_48_n308) );
  FA_X1 mult_48_U140 ( .A(mult_48_n311), .B(mult_48_n391), .CI(mult_48_n308), 
        .CO(mult_48_n305), .S(mult_48_n306) );
  HA_X1 mult_48_U139 ( .A(mult_48_n320), .B(mult_48_n378), .CO(mult_48_n303), 
        .S(mult_48_n304) );
  FA_X1 mult_48_U138 ( .A(mult_48_n390), .B(mult_48_n415), .CI(mult_48_n402), 
        .CO(mult_48_n301), .S(mult_48_n302) );
  FA_X1 mult_48_U137 ( .A(mult_48_n307), .B(mult_48_n304), .CI(mult_48_n302), 
        .CO(mult_48_n299), .S(mult_48_n300) );
  FA_X1 mult_48_U136 ( .A(mult_48_n389), .B(mult_48_n365), .CI(mult_48_n414), 
        .CO(mult_48_n297), .S(mult_48_n298) );
  FA_X1 mult_48_U135 ( .A(mult_48_n377), .B(mult_48_n401), .CI(mult_48_n303), 
        .CO(mult_48_n295), .S(mult_48_n296) );
  FA_X1 mult_48_U134 ( .A(mult_48_n298), .B(mult_48_n301), .CI(mult_48_n296), 
        .CO(mult_48_n293), .S(mult_48_n294) );
  HA_X1 mult_48_U133 ( .A(mult_48_n319), .B(mult_48_n364), .CO(mult_48_n291), 
        .S(mult_48_n292) );
  FA_X1 mult_48_U132 ( .A(mult_48_n376), .B(mult_48_n388), .CI(mult_48_n400), 
        .CO(mult_48_n289), .S(mult_48_n290) );
  FA_X1 mult_48_U131 ( .A(mult_48_n292), .B(mult_48_n413), .CI(mult_48_n297), 
        .CO(mult_48_n287), .S(mult_48_n288) );
  FA_X1 mult_48_U130 ( .A(mult_48_n290), .B(mult_48_n295), .CI(mult_48_n288), 
        .CO(mult_48_n285), .S(mult_48_n286) );
  FA_X1 mult_48_U129 ( .A(mult_48_n375), .B(mult_48_n351), .CI(mult_48_n412), 
        .CO(mult_48_n283), .S(mult_48_n284) );
  FA_X1 mult_48_U128 ( .A(mult_48_n363), .B(mult_48_n399), .CI(mult_48_n387), 
        .CO(mult_48_n281), .S(mult_48_n282) );
  FA_X1 mult_48_U127 ( .A(mult_48_n289), .B(mult_48_n291), .CI(mult_48_n284), 
        .CO(mult_48_n279), .S(mult_48_n280) );
  FA_X1 mult_48_U126 ( .A(mult_48_n287), .B(mult_48_n282), .CI(mult_48_n280), 
        .CO(mult_48_n277), .S(mult_48_n278) );
  HA_X1 mult_48_U125 ( .A(mult_48_n318), .B(mult_48_n350), .CO(mult_48_n275), 
        .S(mult_48_n276) );
  FA_X1 mult_48_U124 ( .A(mult_48_n362), .B(mult_48_n386), .CI(mult_48_n411), 
        .CO(mult_48_n273), .S(mult_48_n274) );
  FA_X1 mult_48_U123 ( .A(mult_48_n374), .B(mult_48_n398), .CI(mult_48_n276), 
        .CO(mult_48_n271), .S(mult_48_n272) );
  FA_X1 mult_48_U122 ( .A(mult_48_n281), .B(mult_48_n283), .CI(mult_48_n274), 
        .CO(mult_48_n269), .S(mult_48_n270) );
  FA_X1 mult_48_U121 ( .A(mult_48_n279), .B(mult_48_n272), .CI(mult_48_n270), 
        .CO(mult_48_n267), .S(mult_48_n268) );
  FA_X1 mult_48_U120 ( .A(mult_48_n361), .B(mult_48_n337), .CI(mult_48_n410), 
        .CO(mult_48_n265), .S(mult_48_n266) );
  FA_X1 mult_48_U109 ( .A(mult_48_n349), .B(mult_48_n397), .CI(mult_48_n373), 
        .CO(mult_48_n263), .S(mult_48_n264) );
  FA_X1 mult_48_U108 ( .A(mult_48_n275), .B(mult_48_n385), .CI(mult_48_n273), 
        .CO(mult_48_n261), .S(mult_48_n262) );
  FA_X1 mult_48_U107 ( .A(mult_48_n264), .B(mult_48_n266), .CI(mult_48_n271), 
        .CO(mult_48_n259), .S(mult_48_n260) );
  FA_X1 mult_48_U106 ( .A(mult_48_n262), .B(mult_48_n269), .CI(mult_48_n260), 
        .CO(mult_48_n257), .S(mult_48_n258) );
  HA_X1 mult_48_U105 ( .A(mult_48_n317), .B(mult_48_n336), .CO(mult_48_n255), 
        .S(mult_48_n256) );
  FA_X1 mult_48_U104 ( .A(mult_48_n409), .B(mult_48_n372), .CI(mult_48_n396), 
        .CO(mult_48_n253), .S(mult_48_n254) );
  FA_X1 mult_48_U103 ( .A(mult_48_n348), .B(mult_48_n384), .CI(mult_48_n360), 
        .CO(mult_48_n251), .S(mult_48_n252) );
  FA_X1 mult_48_U102 ( .A(mult_48_n265), .B(mult_48_n256), .CI(mult_48_n263), 
        .CO(mult_48_n249), .S(mult_48_n250) );
  FA_X1 mult_48_U101 ( .A(mult_48_n254), .B(mult_48_n252), .CI(mult_48_n261), 
        .CO(mult_48_n247), .S(mult_48_n248) );
  FA_X1 mult_48_U100 ( .A(mult_48_n259), .B(mult_48_n250), .CI(mult_48_n248), 
        .CO(mult_48_n245), .S(mult_48_n246) );
  FA_X1 mult_48_U97 ( .A(mult_48_n395), .B(mult_48_n359), .CI(mult_48_n408), 
        .CO(mult_48_n241), .S(mult_48_n242) );
  FA_X1 mult_48_U96 ( .A(mult_48_n335), .B(mult_48_n371), .CI(mult_48_n255), 
        .CO(mult_48_n239), .S(mult_48_n240) );
  FA_X1 mult_48_U95 ( .A(mult_48_n253), .B(mult_48_n244), .CI(mult_48_n251), 
        .CO(mult_48_n237), .S(mult_48_n238) );
  FA_X1 mult_48_U94 ( .A(mult_48_n240), .B(mult_48_n242), .CI(mult_48_n249), 
        .CO(mult_48_n235), .S(mult_48_n236) );
  FA_X1 mult_48_U93 ( .A(mult_48_n247), .B(mult_48_n238), .CI(mult_48_n236), 
        .CO(mult_48_n233), .S(mult_48_n234) );
  FA_X1 mult_48_U91 ( .A(mult_48_n382), .B(mult_48_n346), .CI(mult_48_n232), 
        .CO(mult_48_n229), .S(mult_48_n230) );
  FA_X1 mult_48_U90 ( .A(mult_48_n334), .B(mult_48_n370), .CI(mult_48_n358), 
        .CO(mult_48_n227), .S(mult_48_n228) );
  FA_X1 mult_48_U89 ( .A(mult_48_n241), .B(mult_48_n243), .CI(mult_48_n239), 
        .CO(mult_48_n225), .S(mult_48_n226) );
  FA_X1 mult_48_U88 ( .A(mult_48_n230), .B(mult_48_n228), .CI(mult_48_n237), 
        .CO(mult_48_n223), .S(mult_48_n224) );
  FA_X1 mult_48_U87 ( .A(mult_48_n235), .B(mult_48_n226), .CI(mult_48_n224), 
        .CO(mult_48_n221), .S(mult_48_n222) );
  FA_X1 mult_48_U86 ( .A(mult_48_n231), .B(mult_48_n333), .CI(mult_48_n394), 
        .CO(mult_48_n219), .S(mult_48_n220) );
  FA_X1 mult_48_U85 ( .A(mult_48_n345), .B(mult_48_n381), .CI(mult_48_n357), 
        .CO(mult_48_n217), .S(mult_48_n218) );
  FA_X1 mult_48_U84 ( .A(mult_48_n229), .B(mult_48_n369), .CI(mult_48_n227), 
        .CO(mult_48_n215), .S(mult_48_n216) );
  FA_X1 mult_48_U83 ( .A(mult_48_n220), .B(mult_48_n218), .CI(mult_48_n225), 
        .CO(mult_48_n213), .S(mult_48_n214) );
  FA_X1 mult_48_U82 ( .A(mult_48_n223), .B(mult_48_n216), .CI(mult_48_n214), 
        .CO(mult_48_n211), .S(mult_48_n212) );
  FA_X1 mult_48_U80 ( .A(mult_48_n368), .B(mult_48_n344), .CI(mult_48_n210), 
        .CO(mult_48_n207), .S(mult_48_n208) );
  FA_X1 mult_48_U79 ( .A(mult_48_n332), .B(mult_48_n356), .CI(mult_48_n219), 
        .CO(mult_48_n205), .S(mult_48_n206) );
  FA_X1 mult_48_U78 ( .A(mult_48_n208), .B(mult_48_n217), .CI(mult_48_n215), 
        .CO(mult_48_n203), .S(mult_48_n204) );
  FA_X1 mult_48_U77 ( .A(mult_48_n213), .B(mult_48_n206), .CI(mult_48_n204), 
        .CO(mult_48_n201), .S(mult_48_n202) );
  FA_X1 mult_48_U76 ( .A(mult_48_n209), .B(mult_48_n331), .CI(mult_48_n380), 
        .CO(mult_48_n199), .S(mult_48_n200) );
  FA_X1 mult_48_U75 ( .A(mult_48_n355), .B(mult_48_n343), .CI(mult_48_n367), 
        .CO(mult_48_n197), .S(mult_48_n198) );
  FA_X1 mult_48_U74 ( .A(mult_48_n198), .B(mult_48_n207), .CI(mult_48_n200), 
        .CO(mult_48_n195), .S(mult_48_n196) );
  FA_X1 mult_48_U73 ( .A(mult_48_n203), .B(mult_48_n205), .CI(mult_48_n196), 
        .CO(mult_48_n193), .S(mult_48_n194) );
  FA_X1 mult_48_U71 ( .A(mult_48_n330), .B(mult_48_n342), .CI(mult_48_n192), 
        .CO(mult_48_n189), .S(mult_48_n190) );
  FA_X1 mult_48_U70 ( .A(mult_48_n199), .B(mult_48_n354), .CI(mult_48_n197), 
        .CO(mult_48_n187), .S(mult_48_n188) );
  FA_X1 mult_48_U69 ( .A(mult_48_n188), .B(mult_48_n190), .CI(mult_48_n195), 
        .CO(mult_48_n185), .S(mult_48_n186) );
  FA_X1 mult_48_U68 ( .A(mult_48_n191), .B(mult_48_n329), .CI(mult_48_n366), 
        .CO(mult_48_n183), .S(mult_48_n184) );
  FA_X1 mult_48_U67 ( .A(mult_48_n341), .B(mult_48_n353), .CI(mult_48_n189), 
        .CO(mult_48_n181), .S(mult_48_n182) );
  FA_X1 mult_48_U66 ( .A(mult_48_n187), .B(mult_48_n184), .CI(mult_48_n182), 
        .CO(mult_48_n179), .S(mult_48_n180) );
  FA_X1 mult_48_U64 ( .A(mult_48_n328), .B(mult_48_n340), .CI(mult_48_n178), 
        .CO(mult_48_n175), .S(mult_48_n176) );
  FA_X1 mult_48_U63 ( .A(mult_48_n176), .B(mult_48_n183), .CI(mult_48_n181), 
        .CO(mult_48_n173), .S(mult_48_n174) );
  FA_X1 mult_48_U62 ( .A(mult_48_n327), .B(mult_48_n177), .CI(mult_48_n352), 
        .CO(mult_48_n171), .S(mult_48_n172) );
  FA_X1 mult_48_U61 ( .A(mult_48_n175), .B(mult_48_n339), .CI(mult_48_n172), 
        .CO(mult_48_n169), .S(mult_48_n170) );
  FA_X1 mult_48_U59 ( .A(mult_48_n168), .B(mult_48_n326), .CI(mult_48_n171), 
        .CO(mult_48_n165), .S(mult_48_n166) );
  FA_X1 mult_48_U58 ( .A(mult_48_n325), .B(mult_48_n167), .CI(mult_48_n338), 
        .CO(mult_48_n163), .S(mult_48_n164) );
  FA_X1 mult_48_U44 ( .A(mult_48_n246), .B(mult_48_n257), .CI(mult_48_n149), 
        .CO(mult_48_n148), .S(temp2_13_) );
  FA_X1 mult_48_U43 ( .A(mult_48_n234), .B(mult_48_n245), .CI(mult_48_n148), 
        .CO(mult_48_n147), .S(temp2_14_) );
  FA_X1 mult_48_U42 ( .A(mult_48_n222), .B(mult_48_n233), .CI(mult_48_n147), 
        .CO(mult_48_n146), .S(temp2_15_) );
  FA_X1 mult_48_U41 ( .A(mult_48_n212), .B(mult_48_n221), .CI(mult_48_n146), 
        .CO(mult_48_n145), .S(temp2_16_) );
  FA_X1 mult_48_U40 ( .A(mult_48_n202), .B(mult_48_n211), .CI(mult_48_n145), 
        .CO(mult_48_n144), .S(temp2_17_) );
  FA_X1 mult_48_U39 ( .A(mult_48_n194), .B(mult_48_n201), .CI(mult_48_n144), 
        .CO(mult_48_n143), .S(temp2_18_) );
  FA_X1 mult_48_U38 ( .A(mult_48_n186), .B(mult_48_n193), .CI(mult_48_n143), 
        .CO(mult_48_n142), .S(temp2_19_) );
  FA_X1 mult_48_U37 ( .A(mult_48_n180), .B(mult_48_n185), .CI(mult_48_n142), 
        .CO(mult_48_n141), .S(temp2_20_) );
  FA_X1 mult_48_U30 ( .A(mult_48_n174), .B(mult_48_n179), .CI(mult_48_n141), 
        .CO(mult_48_n140), .S(temp2_21_) );
  FA_X1 mult_48_U20 ( .A(mult_48_n170), .B(mult_48_n173), .CI(mult_48_n140), 
        .CO(mult_48_n139), .S(temp2_22_) );
  FA_X1 mult_48_U10 ( .A(mult_48_n166), .B(mult_48_n169), .CI(mult_48_n139), 
        .CO(mult_48_n138), .S(temp2_23_) );
  FA_X1 mult_48_U9 ( .A(mult_48_n165), .B(mult_48_n164), .CI(mult_48_n138), 
        .CO(mult_48_n137), .S(temp2_24_) );
  FA_X1 mult_48_U8 ( .A(mult_48_n163), .B(mult_48_n162), .CI(mult_48_n137), 
        .CO(mult_48_n136), .S(temp2_25_) );
  INV_X1 sub_1_root_add_0_root_add_58_U16 ( .A(temp1_13_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_0_) );
  INV_X1 sub_1_root_add_0_root_add_58_U15 ( .A(temp1_23_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_10_) );
  INV_X1 sub_1_root_add_0_root_add_58_U14 ( .A(temp1_24_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_11_) );
  INV_X1 sub_1_root_add_0_root_add_58_U13 ( .A(temp1_25_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_12_) );
  INV_X1 sub_1_root_add_0_root_add_58_U12 ( .A(temp1_26_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_13_) );
  INV_X1 sub_1_root_add_0_root_add_58_U11 ( .A(temp1_14_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_1_) );
  INV_X1 sub_1_root_add_0_root_add_58_U10 ( .A(temp1_15_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_2_) );
  INV_X1 sub_1_root_add_0_root_add_58_U9 ( .A(temp1_16_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_3_) );
  INV_X1 sub_1_root_add_0_root_add_58_U8 ( .A(temp1_17_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_4_) );
  INV_X1 sub_1_root_add_0_root_add_58_U7 ( .A(temp1_18_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_5_) );
  INV_X1 sub_1_root_add_0_root_add_58_U6 ( .A(temp1_19_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_6_) );
  INV_X1 sub_1_root_add_0_root_add_58_U5 ( .A(temp1_20_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_7_) );
  INV_X1 sub_1_root_add_0_root_add_58_U4 ( .A(temp1_21_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_8_) );
  INV_X1 sub_1_root_add_0_root_add_58_U3 ( .A(temp1_22_), .ZN(
        sub_1_root_add_0_root_add_58_B_not_9_) );
  XNOR2_X1 sub_1_root_add_0_root_add_58_U2 ( .A(fb_0_), .B(
        sub_1_root_add_0_root_add_58_B_not_0_), .ZN(N0) );
  OR2_X1 sub_1_root_add_0_root_add_58_U1 ( .A1(
        sub_1_root_add_0_root_add_58_B_not_0_), .A2(fb_0_), .ZN(
        sub_1_root_add_0_root_add_58_carry_1_) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_1 ( .A(fb_1_), .B(
        sub_1_root_add_0_root_add_58_B_not_1_), .CI(
        sub_1_root_add_0_root_add_58_carry_1_), .CO(
        sub_1_root_add_0_root_add_58_carry_2_), .S(N1) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_2 ( .A(fb_2_), .B(
        sub_1_root_add_0_root_add_58_B_not_2_), .CI(
        sub_1_root_add_0_root_add_58_carry_2_), .CO(
        sub_1_root_add_0_root_add_58_carry_3_), .S(N2) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_3 ( .A(fb_3_), .B(
        sub_1_root_add_0_root_add_58_B_not_3_), .CI(
        sub_1_root_add_0_root_add_58_carry_3_), .CO(
        sub_1_root_add_0_root_add_58_carry_4_), .S(N3) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_4 ( .A(fb_4_), .B(
        sub_1_root_add_0_root_add_58_B_not_4_), .CI(
        sub_1_root_add_0_root_add_58_carry_4_), .CO(
        sub_1_root_add_0_root_add_58_carry_5_), .S(N4) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_5 ( .A(fb_5_), .B(
        sub_1_root_add_0_root_add_58_B_not_5_), .CI(
        sub_1_root_add_0_root_add_58_carry_5_), .CO(
        sub_1_root_add_0_root_add_58_carry_6_), .S(N5) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_6 ( .A(fb_6_), .B(
        sub_1_root_add_0_root_add_58_B_not_6_), .CI(
        sub_1_root_add_0_root_add_58_carry_6_), .CO(
        sub_1_root_add_0_root_add_58_carry_7_), .S(N6) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_7 ( .A(fb_7_), .B(
        sub_1_root_add_0_root_add_58_B_not_7_), .CI(
        sub_1_root_add_0_root_add_58_carry_7_), .CO(
        sub_1_root_add_0_root_add_58_carry_8_), .S(N7) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_8 ( .A(fb_8_), .B(
        sub_1_root_add_0_root_add_58_B_not_8_), .CI(
        sub_1_root_add_0_root_add_58_carry_8_), .CO(
        sub_1_root_add_0_root_add_58_carry_9_), .S(N8) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_9 ( .A(fb_9_), .B(
        sub_1_root_add_0_root_add_58_B_not_9_), .CI(
        sub_1_root_add_0_root_add_58_carry_9_), .CO(
        sub_1_root_add_0_root_add_58_carry_10_), .S(N9) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_10 ( .A(fb_10_), .B(
        sub_1_root_add_0_root_add_58_B_not_10_), .CI(
        sub_1_root_add_0_root_add_58_carry_10_), .CO(
        sub_1_root_add_0_root_add_58_carry_11_), .S(N10) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_11 ( .A(fb_11_), .B(
        sub_1_root_add_0_root_add_58_B_not_11_), .CI(
        sub_1_root_add_0_root_add_58_carry_11_), .CO(
        sub_1_root_add_0_root_add_58_carry_12_), .S(N11) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_12 ( .A(fb_12_), .B(
        sub_1_root_add_0_root_add_58_B_not_12_), .CI(
        sub_1_root_add_0_root_add_58_carry_12_), .CO(
        sub_1_root_add_0_root_add_58_carry_13_), .S(N12) );
  FA_X1 sub_1_root_add_0_root_add_58_U2_13 ( .A(fb_13_), .B(
        sub_1_root_add_0_root_add_58_B_not_13_), .CI(
        sub_1_root_add_0_root_add_58_carry_13_), .S(N13) );
  INV_X1 sub_0_root_add_0_root_add_58_U16 ( .A(temp2_13_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_0_) );
  INV_X1 sub_0_root_add_0_root_add_58_U15 ( .A(temp2_23_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_10_) );
  INV_X1 sub_0_root_add_0_root_add_58_U14 ( .A(temp2_24_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_11_) );
  INV_X1 sub_0_root_add_0_root_add_58_U13 ( .A(temp2_25_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_12_) );
  INV_X1 sub_0_root_add_0_root_add_58_U12 ( .A(temp2_26_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_13_) );
  INV_X1 sub_0_root_add_0_root_add_58_U11 ( .A(temp2_14_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_1_) );
  INV_X1 sub_0_root_add_0_root_add_58_U10 ( .A(temp2_15_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_2_) );
  INV_X1 sub_0_root_add_0_root_add_58_U9 ( .A(temp2_16_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_3_) );
  INV_X1 sub_0_root_add_0_root_add_58_U8 ( .A(temp2_17_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_4_) );
  INV_X1 sub_0_root_add_0_root_add_58_U7 ( .A(temp2_18_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_5_) );
  INV_X1 sub_0_root_add_0_root_add_58_U6 ( .A(temp2_19_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_6_) );
  INV_X1 sub_0_root_add_0_root_add_58_U5 ( .A(temp2_20_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_7_) );
  INV_X1 sub_0_root_add_0_root_add_58_U4 ( .A(temp2_21_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_8_) );
  INV_X1 sub_0_root_add_0_root_add_58_U3 ( .A(temp2_22_), .ZN(
        sub_0_root_add_0_root_add_58_B_not_9_) );
  XNOR2_X1 sub_0_root_add_0_root_add_58_U2 ( .A(N0), .B(
        sub_0_root_add_0_root_add_58_B_not_0_), .ZN(w[0]) );
  OR2_X1 sub_0_root_add_0_root_add_58_U1 ( .A1(
        sub_0_root_add_0_root_add_58_B_not_0_), .A2(N0), .ZN(
        sub_0_root_add_0_root_add_58_carry_1_) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_1 ( .A(N1), .B(
        sub_0_root_add_0_root_add_58_B_not_1_), .CI(
        sub_0_root_add_0_root_add_58_carry_1_), .CO(
        sub_0_root_add_0_root_add_58_carry_2_), .S(w[1]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_2 ( .A(N2), .B(
        sub_0_root_add_0_root_add_58_B_not_2_), .CI(
        sub_0_root_add_0_root_add_58_carry_2_), .CO(
        sub_0_root_add_0_root_add_58_carry_3_), .S(w[2]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_3 ( .A(N3), .B(
        sub_0_root_add_0_root_add_58_B_not_3_), .CI(
        sub_0_root_add_0_root_add_58_carry_3_), .CO(
        sub_0_root_add_0_root_add_58_carry_4_), .S(w[3]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_4 ( .A(N4), .B(
        sub_0_root_add_0_root_add_58_B_not_4_), .CI(
        sub_0_root_add_0_root_add_58_carry_4_), .CO(
        sub_0_root_add_0_root_add_58_carry_5_), .S(w[4]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_5 ( .A(N5), .B(
        sub_0_root_add_0_root_add_58_B_not_5_), .CI(
        sub_0_root_add_0_root_add_58_carry_5_), .CO(
        sub_0_root_add_0_root_add_58_carry_6_), .S(w[5]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_6 ( .A(N6), .B(
        sub_0_root_add_0_root_add_58_B_not_6_), .CI(
        sub_0_root_add_0_root_add_58_carry_6_), .CO(
        sub_0_root_add_0_root_add_58_carry_7_), .S(w[6]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_7 ( .A(N7), .B(
        sub_0_root_add_0_root_add_58_B_not_7_), .CI(
        sub_0_root_add_0_root_add_58_carry_7_), .CO(
        sub_0_root_add_0_root_add_58_carry_8_), .S(w[7]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_8 ( .A(N8), .B(
        sub_0_root_add_0_root_add_58_B_not_8_), .CI(
        sub_0_root_add_0_root_add_58_carry_8_), .CO(
        sub_0_root_add_0_root_add_58_carry_9_), .S(w[8]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_9 ( .A(N9), .B(
        sub_0_root_add_0_root_add_58_B_not_9_), .CI(
        sub_0_root_add_0_root_add_58_carry_9_), .CO(
        sub_0_root_add_0_root_add_58_carry_10_), .S(w[9]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_10 ( .A(N10), .B(
        sub_0_root_add_0_root_add_58_B_not_10_), .CI(
        sub_0_root_add_0_root_add_58_carry_10_), .CO(
        sub_0_root_add_0_root_add_58_carry_11_), .S(w[10]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_11 ( .A(N11), .B(
        sub_0_root_add_0_root_add_58_B_not_11_), .CI(
        sub_0_root_add_0_root_add_58_carry_11_), .CO(
        sub_0_root_add_0_root_add_58_carry_12_), .S(w[11]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_12 ( .A(N12), .B(
        sub_0_root_add_0_root_add_58_B_not_12_), .CI(
        sub_0_root_add_0_root_add_58_carry_12_), .CO(
        sub_0_root_add_0_root_add_58_carry_13_), .S(w[12]) );
  FA_X1 sub_0_root_add_0_root_add_58_U2_13 ( .A(N13), .B(
        sub_0_root_add_0_root_add_58_B_not_13_), .CI(
        sub_0_root_add_0_root_add_58_carry_13_), .S(w[13]) );
endmodule

