
module IIR_ADV ( CLK, RST_n, VIN, DIN, B0, B1, B2, B3, A1, A2, VOUT, DOUT );
  input [13:0] DIN;
  input [13:0] B0;
  input [13:0] B1;
  input [13:0] B2;
  input [13:0] B3;
  input [13:0] A1;
  input [13:0] A2;
  output [13:0] DOUT;
  input CLK, RST_n, VIN;
  output VOUT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, REGISTER1_n47, REGISTER1_n46, REGISTER1_n45,
         REGISTER1_n44, REGISTER1_n43, REGISTER1_n42, REGISTER1_n41,
         REGISTER1_n40, REGISTER1_n39, REGISTER1_n38, REGISTER1_n37,
         REGISTER1_n36, REGISTER1_n35, REGISTER1_n34, REGISTER1_n33,
         REGISTER1_n32, REGISTER1_n31, REGISTER1_n30, REGISTER1_n29,
         REGISTER1_n28, REGISTER1_n27, REGISTER1_n26, REGISTER1_n25,
         REGISTER1_n24, REGISTER1_n23, REGISTER1_n22, REGISTER1_n21,
         REGISTER1_n20, REGISTER1_n19, REGISTER1_n18, REGISTER1_n17,
         REGISTER1_n16, REGISTER1_n15, REGISTER1_n14, REGISTER1_n13,
         REGISTER1_n12, REGISTER1_n11, REGISTER1_n10, REGISTER1_n9,
         REGISTER1_n8, REGISTER1_n7, REGISTER1_n6, REGISTER1_n5, REGISTER1_n4,
         REGISTER1_n3, REGISTER1_n2, REGISTER1_n1, p6_mult_21_n805,
         p6_mult_21_n804, p6_mult_21_n803, p6_mult_21_n802, p6_mult_21_n801,
         p6_mult_21_n800, p6_mult_21_n799, p6_mult_21_n798, p6_mult_21_n797,
         p6_mult_21_n796, p6_mult_21_n795, p6_mult_21_n794, p6_mult_21_n793,
         p6_mult_21_n792, p6_mult_21_n791, p6_mult_21_n790, p6_mult_21_n789,
         p6_mult_21_n788, p6_mult_21_n787, p6_mult_21_n786, p6_mult_21_n785,
         p6_mult_21_n784, p6_mult_21_n783, p6_mult_21_n782, p6_mult_21_n781,
         p6_mult_21_n780, p6_mult_21_n779, p6_mult_21_n778, p6_mult_21_n777,
         p6_mult_21_n776, p6_mult_21_n775, p6_mult_21_n774, p6_mult_21_n773,
         p6_mult_21_n772, p6_mult_21_n771, p6_mult_21_n770, p6_mult_21_n769,
         p6_mult_21_n768, p6_mult_21_n767, p6_mult_21_n766, p6_mult_21_n765,
         p6_mult_21_n764, p6_mult_21_n763, p6_mult_21_n762, p6_mult_21_n761,
         p6_mult_21_n760, p6_mult_21_n759, p6_mult_21_n758, p6_mult_21_n757,
         p6_mult_21_n756, p6_mult_21_n755, p6_mult_21_n754, p6_mult_21_n753,
         p6_mult_21_n752, p6_mult_21_n751, p6_mult_21_n750, p6_mult_21_n749,
         p6_mult_21_n748, p6_mult_21_n747, p6_mult_21_n746, p6_mult_21_n745,
         p6_mult_21_n744, p6_mult_21_n743, p6_mult_21_n742, p6_mult_21_n741,
         p6_mult_21_n740, p6_mult_21_n739, p6_mult_21_n738, p6_mult_21_n737,
         p6_mult_21_n736, p6_mult_21_n735, p6_mult_21_n734, p6_mult_21_n733,
         p6_mult_21_n732, p6_mult_21_n731, p6_mult_21_n730, p6_mult_21_n729,
         p6_mult_21_n728, p6_mult_21_n727, p6_mult_21_n726, p6_mult_21_n725,
         p6_mult_21_n724, p6_mult_21_n723, p6_mult_21_n722, p6_mult_21_n721,
         p6_mult_21_n720, p6_mult_21_n719, p6_mult_21_n718, p6_mult_21_n717,
         p6_mult_21_n716, p6_mult_21_n715, p6_mult_21_n714, p6_mult_21_n713,
         p6_mult_21_n712, p6_mult_21_n711, p6_mult_21_n710, p6_mult_21_n709,
         p6_mult_21_n708, p6_mult_21_n707, p6_mult_21_n706, p6_mult_21_n705,
         p6_mult_21_n704, p6_mult_21_n703, p6_mult_21_n702, p6_mult_21_n701,
         p6_mult_21_n700, p6_mult_21_n699, p6_mult_21_n698, p6_mult_21_n697,
         p6_mult_21_n696, p6_mult_21_n695, p6_mult_21_n694, p6_mult_21_n693,
         p6_mult_21_n692, p6_mult_21_n691, p6_mult_21_n690, p6_mult_21_n689,
         p6_mult_21_n688, p6_mult_21_n687, p6_mult_21_n686, p6_mult_21_n685,
         p6_mult_21_n684, p6_mult_21_n683, p6_mult_21_n682, p6_mult_21_n681,
         p6_mult_21_n680, p6_mult_21_n679, p6_mult_21_n678, p6_mult_21_n677,
         p6_mult_21_n676, p6_mult_21_n675, p6_mult_21_n674, p6_mult_21_n673,
         p6_mult_21_n672, p6_mult_21_n671, p6_mult_21_n670, p6_mult_21_n669,
         p6_mult_21_n668, p6_mult_21_n667, p6_mult_21_n666, p6_mult_21_n665,
         p6_mult_21_n664, p6_mult_21_n663, p6_mult_21_n662, p6_mult_21_n661,
         p6_mult_21_n660, p6_mult_21_n659, p6_mult_21_n658, p6_mult_21_n657,
         p6_mult_21_n656, p6_mult_21_n655, p6_mult_21_n654, p6_mult_21_n653,
         p6_mult_21_n652, p6_mult_21_n651, p6_mult_21_n650, p6_mult_21_n649,
         p6_mult_21_n648, p6_mult_21_n647, p6_mult_21_n646, p6_mult_21_n645,
         p6_mult_21_n644, p6_mult_21_n643, p6_mult_21_n642, p6_mult_21_n641,
         p6_mult_21_n640, p6_mult_21_n639, p6_mult_21_n638, p6_mult_21_n637,
         p6_mult_21_n636, p6_mult_21_n635, p6_mult_21_n419, p6_mult_21_n418,
         p6_mult_21_n417, p6_mult_21_n416, p6_mult_21_n415, p6_mult_21_n414,
         p6_mult_21_n413, p6_mult_21_n412, p6_mult_21_n411, p6_mult_21_n410,
         p6_mult_21_n409, p6_mult_21_n408, p6_mult_21_n406, p6_mult_21_n405,
         p6_mult_21_n404, p6_mult_21_n403, p6_mult_21_n402, p6_mult_21_n401,
         p6_mult_21_n400, p6_mult_21_n399, p6_mult_21_n398, p6_mult_21_n397,
         p6_mult_21_n396, p6_mult_21_n395, p6_mult_21_n394, p6_mult_21_n393,
         p6_mult_21_n392, p6_mult_21_n391, p6_mult_21_n390, p6_mult_21_n389,
         p6_mult_21_n388, p6_mult_21_n387, p6_mult_21_n386, p6_mult_21_n385,
         p6_mult_21_n384, p6_mult_21_n382, p6_mult_21_n381, p6_mult_21_n380,
         p6_mult_21_n379, p6_mult_21_n378, p6_mult_21_n377, p6_mult_21_n376,
         p6_mult_21_n375, p6_mult_21_n374, p6_mult_21_n373, p6_mult_21_n372,
         p6_mult_21_n371, p6_mult_21_n370, p6_mult_21_n369, p6_mult_21_n368,
         p6_mult_21_n367, p6_mult_21_n366, p6_mult_21_n365, p6_mult_21_n364,
         p6_mult_21_n363, p6_mult_21_n362, p6_mult_21_n361, p6_mult_21_n360,
         p6_mult_21_n359, p6_mult_21_n358, p6_mult_21_n357, p6_mult_21_n356,
         p6_mult_21_n355, p6_mult_21_n354, p6_mult_21_n353, p6_mult_21_n352,
         p6_mult_21_n351, p6_mult_21_n350, p6_mult_21_n349, p6_mult_21_n348,
         p6_mult_21_n346, p6_mult_21_n345, p6_mult_21_n344, p6_mult_21_n343,
         p6_mult_21_n342, p6_mult_21_n341, p6_mult_21_n340, p6_mult_21_n339,
         p6_mult_21_n338, p6_mult_21_n337, p6_mult_21_n336, p6_mult_21_n335,
         p6_mult_21_n334, p6_mult_21_n333, p6_mult_21_n332, p6_mult_21_n331,
         p6_mult_21_n330, p6_mult_21_n329, p6_mult_21_n328, p6_mult_21_n327,
         p6_mult_21_n326, p6_mult_21_n325, p6_mult_21_n321, p6_mult_21_n320,
         p6_mult_21_n319, p6_mult_21_n318, p6_mult_21_n317, p6_mult_21_n316,
         p6_mult_21_n315, p6_mult_21_n314, p6_mult_21_n313, p6_mult_21_n312,
         p6_mult_21_n311, p6_mult_21_n310, p6_mult_21_n309, p6_mult_21_n308,
         p6_mult_21_n307, p6_mult_21_n306, p6_mult_21_n305, p6_mult_21_n304,
         p6_mult_21_n303, p6_mult_21_n302, p6_mult_21_n301, p6_mult_21_n300,
         p6_mult_21_n299, p6_mult_21_n298, p6_mult_21_n297, p6_mult_21_n296,
         p6_mult_21_n295, p6_mult_21_n294, p6_mult_21_n293, p6_mult_21_n292,
         p6_mult_21_n291, p6_mult_21_n290, p6_mult_21_n289, p6_mult_21_n288,
         p6_mult_21_n287, p6_mult_21_n286, p6_mult_21_n285, p6_mult_21_n284,
         p6_mult_21_n283, p6_mult_21_n282, p6_mult_21_n281, p6_mult_21_n280,
         p6_mult_21_n279, p6_mult_21_n278, p6_mult_21_n277, p6_mult_21_n276,
         p6_mult_21_n275, p6_mult_21_n274, p6_mult_21_n273, p6_mult_21_n272,
         p6_mult_21_n271, p6_mult_21_n270, p6_mult_21_n269, p6_mult_21_n268,
         p6_mult_21_n267, p6_mult_21_n266, p6_mult_21_n265, p6_mult_21_n264,
         p6_mult_21_n263, p6_mult_21_n262, p6_mult_21_n261, p6_mult_21_n260,
         p6_mult_21_n259, p6_mult_21_n258, p6_mult_21_n257, p6_mult_21_n256,
         p6_mult_21_n255, p6_mult_21_n254, p6_mult_21_n253, p6_mult_21_n252,
         p6_mult_21_n251, p6_mult_21_n250, p6_mult_21_n249, p6_mult_21_n248,
         p6_mult_21_n247, p6_mult_21_n246, p6_mult_21_n245, p6_mult_21_n244,
         p6_mult_21_n243, p6_mult_21_n242, p6_mult_21_n241, p6_mult_21_n240,
         p6_mult_21_n239, p6_mult_21_n238, p6_mult_21_n237, p6_mult_21_n236,
         p6_mult_21_n235, p6_mult_21_n234, p6_mult_21_n233, p6_mult_21_n232,
         p6_mult_21_n231, p6_mult_21_n230, p6_mult_21_n229, p6_mult_21_n228,
         p6_mult_21_n227, p6_mult_21_n226, p6_mult_21_n225, p6_mult_21_n224,
         p6_mult_21_n223, p6_mult_21_n222, p6_mult_21_n221, p6_mult_21_n220,
         p6_mult_21_n219, p6_mult_21_n218, p6_mult_21_n217, p6_mult_21_n216,
         p6_mult_21_n215, p6_mult_21_n214, p6_mult_21_n213, p6_mult_21_n212,
         p6_mult_21_n211, p6_mult_21_n210, p6_mult_21_n209, p6_mult_21_n208,
         p6_mult_21_n207, p6_mult_21_n206, p6_mult_21_n205, p6_mult_21_n204,
         p6_mult_21_n203, p6_mult_21_n202, p6_mult_21_n201, p6_mult_21_n200,
         p6_mult_21_n199, p6_mult_21_n198, p6_mult_21_n197, p6_mult_21_n196,
         p6_mult_21_n195, p6_mult_21_n194, p6_mult_21_n193, p6_mult_21_n192,
         p6_mult_21_n191, p6_mult_21_n190, p6_mult_21_n189, p6_mult_21_n188,
         p6_mult_21_n187, p6_mult_21_n186, p6_mult_21_n185, p6_mult_21_n184,
         p6_mult_21_n183, p6_mult_21_n182, p6_mult_21_n181, p6_mult_21_n180,
         p6_mult_21_n179, p6_mult_21_n178, p6_mult_21_n177, p6_mult_21_n176,
         p6_mult_21_n175, p6_mult_21_n174, p6_mult_21_n173, p6_mult_21_n172,
         p6_mult_21_n171, p6_mult_21_n170, p6_mult_21_n169, p6_mult_21_n168,
         p6_mult_21_n167, p6_mult_21_n166, p6_mult_21_n165, p6_mult_21_n164,
         p6_mult_21_n163, p6_mult_21_n162, p6_mult_21_n149, p6_mult_21_n148,
         p6_mult_21_n147, p6_mult_21_n146, p6_mult_21_n145, p6_mult_21_n144,
         p6_mult_21_n143, p6_mult_21_n142, p6_mult_21_n141, p6_mult_21_n140,
         p6_mult_21_n139, p6_mult_21_n138, p6_mult_21_n137, p6_mult_21_n136,
         REG1_1_n89, REG1_1_n88, REG1_1_n87, REG1_1_n86, REG1_1_n85,
         REG1_1_n84, REG1_1_n83, REG1_1_n82, REG1_1_n81, REG1_1_n80,
         REG1_1_n79, REG1_1_n78, REG1_1_n77, REG1_1_n76, REG1_1_n75,
         REG1_1_n74, REG1_1_n73, REG1_1_n72, REG1_1_n71, REG1_1_n70,
         REG1_1_n69, REG1_1_n68, REG1_1_n67, REG1_1_n66, REG1_1_n65,
         REG1_1_n64, REG1_1_n63, REG1_1_n62, REG1_1_n61, REG1_1_n60,
         REG1_1_n59, REG1_1_n58, REG1_1_n57, REG1_1_n56, REG1_1_n55,
         REG1_1_n54, REG1_1_n53, REG1_1_n52, REG1_1_n51, REG1_1_n50,
         REG1_1_n49, REG1_1_n48, REG1_1_n47, REG1_1_n46, REG1_1_n45,
         REG1_1_n44, REG1_1_n43, REGISTER2_n89, REGISTER2_n88, REGISTER2_n87,
         REGISTER2_n86, REGISTER2_n85, REGISTER2_n84, REGISTER2_n83,
         REGISTER2_n82, REGISTER2_n81, REGISTER2_n80, REGISTER2_n79,
         REGISTER2_n78, REGISTER2_n77, REGISTER2_n76, REGISTER2_n75,
         REGISTER2_n74, REGISTER2_n73, REGISTER2_n72, REGISTER2_n71,
         REGISTER2_n70, REGISTER2_n69, REGISTER2_n68, REGISTER2_n67,
         REGISTER2_n66, REGISTER2_n65, REGISTER2_n64, REGISTER2_n63,
         REGISTER2_n62, REGISTER2_n61, REGISTER2_n60, REGISTER2_n59,
         REGISTER2_n58, REGISTER2_n57, REGISTER2_n56, REGISTER2_n55,
         REGISTER2_n54, REGISTER2_n53, REGISTER2_n52, REGISTER2_n51,
         REGISTER2_n50, REGISTER2_n49, REGISTER2_n48, REGISTER2_n47,
         REGISTER2_n46, REGISTER2_n45, REGISTER2_n44, REGISTER2_n43,
         p7_mult_21_n805, p7_mult_21_n804, p7_mult_21_n803, p7_mult_21_n802,
         p7_mult_21_n801, p7_mult_21_n800, p7_mult_21_n799, p7_mult_21_n798,
         p7_mult_21_n797, p7_mult_21_n796, p7_mult_21_n795, p7_mult_21_n794,
         p7_mult_21_n793, p7_mult_21_n792, p7_mult_21_n791, p7_mult_21_n790,
         p7_mult_21_n789, p7_mult_21_n788, p7_mult_21_n787, p7_mult_21_n786,
         p7_mult_21_n785, p7_mult_21_n784, p7_mult_21_n783, p7_mult_21_n782,
         p7_mult_21_n781, p7_mult_21_n780, p7_mult_21_n779, p7_mult_21_n778,
         p7_mult_21_n777, p7_mult_21_n776, p7_mult_21_n775, p7_mult_21_n774,
         p7_mult_21_n773, p7_mult_21_n772, p7_mult_21_n771, p7_mult_21_n770,
         p7_mult_21_n769, p7_mult_21_n768, p7_mult_21_n767, p7_mult_21_n766,
         p7_mult_21_n765, p7_mult_21_n764, p7_mult_21_n763, p7_mult_21_n762,
         p7_mult_21_n761, p7_mult_21_n760, p7_mult_21_n759, p7_mult_21_n758,
         p7_mult_21_n757, p7_mult_21_n756, p7_mult_21_n755, p7_mult_21_n754,
         p7_mult_21_n753, p7_mult_21_n752, p7_mult_21_n751, p7_mult_21_n750,
         p7_mult_21_n749, p7_mult_21_n748, p7_mult_21_n747, p7_mult_21_n746,
         p7_mult_21_n745, p7_mult_21_n744, p7_mult_21_n743, p7_mult_21_n742,
         p7_mult_21_n741, p7_mult_21_n740, p7_mult_21_n739, p7_mult_21_n738,
         p7_mult_21_n737, p7_mult_21_n736, p7_mult_21_n735, p7_mult_21_n734,
         p7_mult_21_n733, p7_mult_21_n732, p7_mult_21_n731, p7_mult_21_n730,
         p7_mult_21_n729, p7_mult_21_n728, p7_mult_21_n727, p7_mult_21_n726,
         p7_mult_21_n725, p7_mult_21_n724, p7_mult_21_n723, p7_mult_21_n722,
         p7_mult_21_n721, p7_mult_21_n720, p7_mult_21_n719, p7_mult_21_n718,
         p7_mult_21_n717, p7_mult_21_n716, p7_mult_21_n715, p7_mult_21_n714,
         p7_mult_21_n713, p7_mult_21_n712, p7_mult_21_n711, p7_mult_21_n710,
         p7_mult_21_n709, p7_mult_21_n708, p7_mult_21_n707, p7_mult_21_n706,
         p7_mult_21_n705, p7_mult_21_n704, p7_mult_21_n703, p7_mult_21_n702,
         p7_mult_21_n701, p7_mult_21_n700, p7_mult_21_n699, p7_mult_21_n698,
         p7_mult_21_n697, p7_mult_21_n696, p7_mult_21_n695, p7_mult_21_n694,
         p7_mult_21_n693, p7_mult_21_n692, p7_mult_21_n691, p7_mult_21_n690,
         p7_mult_21_n689, p7_mult_21_n688, p7_mult_21_n687, p7_mult_21_n686,
         p7_mult_21_n685, p7_mult_21_n684, p7_mult_21_n683, p7_mult_21_n682,
         p7_mult_21_n681, p7_mult_21_n680, p7_mult_21_n679, p7_mult_21_n678,
         p7_mult_21_n677, p7_mult_21_n676, p7_mult_21_n675, p7_mult_21_n674,
         p7_mult_21_n673, p7_mult_21_n672, p7_mult_21_n671, p7_mult_21_n670,
         p7_mult_21_n669, p7_mult_21_n668, p7_mult_21_n667, p7_mult_21_n666,
         p7_mult_21_n665, p7_mult_21_n664, p7_mult_21_n663, p7_mult_21_n662,
         p7_mult_21_n661, p7_mult_21_n660, p7_mult_21_n659, p7_mult_21_n658,
         p7_mult_21_n657, p7_mult_21_n656, p7_mult_21_n655, p7_mult_21_n654,
         p7_mult_21_n653, p7_mult_21_n652, p7_mult_21_n651, p7_mult_21_n650,
         p7_mult_21_n649, p7_mult_21_n648, p7_mult_21_n647, p7_mult_21_n646,
         p7_mult_21_n645, p7_mult_21_n644, p7_mult_21_n643, p7_mult_21_n642,
         p7_mult_21_n641, p7_mult_21_n640, p7_mult_21_n639, p7_mult_21_n638,
         p7_mult_21_n637, p7_mult_21_n636, p7_mult_21_n635, p7_mult_21_n419,
         p7_mult_21_n418, p7_mult_21_n417, p7_mult_21_n416, p7_mult_21_n415,
         p7_mult_21_n414, p7_mult_21_n413, p7_mult_21_n412, p7_mult_21_n411,
         p7_mult_21_n410, p7_mult_21_n409, p7_mult_21_n408, p7_mult_21_n406,
         p7_mult_21_n405, p7_mult_21_n404, p7_mult_21_n403, p7_mult_21_n402,
         p7_mult_21_n401, p7_mult_21_n400, p7_mult_21_n399, p7_mult_21_n398,
         p7_mult_21_n397, p7_mult_21_n396, p7_mult_21_n395, p7_mult_21_n394,
         p7_mult_21_n393, p7_mult_21_n392, p7_mult_21_n391, p7_mult_21_n390,
         p7_mult_21_n389, p7_mult_21_n388, p7_mult_21_n387, p7_mult_21_n386,
         p7_mult_21_n385, p7_mult_21_n384, p7_mult_21_n382, p7_mult_21_n381,
         p7_mult_21_n380, p7_mult_21_n379, p7_mult_21_n378, p7_mult_21_n377,
         p7_mult_21_n376, p7_mult_21_n375, p7_mult_21_n374, p7_mult_21_n373,
         p7_mult_21_n372, p7_mult_21_n371, p7_mult_21_n370, p7_mult_21_n369,
         p7_mult_21_n368, p7_mult_21_n367, p7_mult_21_n366, p7_mult_21_n365,
         p7_mult_21_n364, p7_mult_21_n363, p7_mult_21_n362, p7_mult_21_n361,
         p7_mult_21_n360, p7_mult_21_n359, p7_mult_21_n358, p7_mult_21_n357,
         p7_mult_21_n356, p7_mult_21_n355, p7_mult_21_n354, p7_mult_21_n353,
         p7_mult_21_n352, p7_mult_21_n351, p7_mult_21_n350, p7_mult_21_n349,
         p7_mult_21_n348, p7_mult_21_n346, p7_mult_21_n345, p7_mult_21_n344,
         p7_mult_21_n343, p7_mult_21_n342, p7_mult_21_n341, p7_mult_21_n340,
         p7_mult_21_n339, p7_mult_21_n338, p7_mult_21_n337, p7_mult_21_n336,
         p7_mult_21_n335, p7_mult_21_n334, p7_mult_21_n333, p7_mult_21_n332,
         p7_mult_21_n331, p7_mult_21_n330, p7_mult_21_n329, p7_mult_21_n328,
         p7_mult_21_n327, p7_mult_21_n326, p7_mult_21_n325, p7_mult_21_n321,
         p7_mult_21_n320, p7_mult_21_n319, p7_mult_21_n318, p7_mult_21_n317,
         p7_mult_21_n316, p7_mult_21_n315, p7_mult_21_n314, p7_mult_21_n313,
         p7_mult_21_n312, p7_mult_21_n311, p7_mult_21_n310, p7_mult_21_n309,
         p7_mult_21_n308, p7_mult_21_n307, p7_mult_21_n306, p7_mult_21_n305,
         p7_mult_21_n304, p7_mult_21_n303, p7_mult_21_n302, p7_mult_21_n301,
         p7_mult_21_n300, p7_mult_21_n299, p7_mult_21_n298, p7_mult_21_n297,
         p7_mult_21_n296, p7_mult_21_n295, p7_mult_21_n294, p7_mult_21_n293,
         p7_mult_21_n292, p7_mult_21_n291, p7_mult_21_n290, p7_mult_21_n289,
         p7_mult_21_n288, p7_mult_21_n287, p7_mult_21_n286, p7_mult_21_n285,
         p7_mult_21_n284, p7_mult_21_n283, p7_mult_21_n282, p7_mult_21_n281,
         p7_mult_21_n280, p7_mult_21_n279, p7_mult_21_n278, p7_mult_21_n277,
         p7_mult_21_n276, p7_mult_21_n275, p7_mult_21_n274, p7_mult_21_n273,
         p7_mult_21_n272, p7_mult_21_n271, p7_mult_21_n270, p7_mult_21_n269,
         p7_mult_21_n268, p7_mult_21_n267, p7_mult_21_n266, p7_mult_21_n265,
         p7_mult_21_n264, p7_mult_21_n263, p7_mult_21_n262, p7_mult_21_n261,
         p7_mult_21_n260, p7_mult_21_n259, p7_mult_21_n258, p7_mult_21_n257,
         p7_mult_21_n256, p7_mult_21_n255, p7_mult_21_n254, p7_mult_21_n253,
         p7_mult_21_n252, p7_mult_21_n251, p7_mult_21_n250, p7_mult_21_n249,
         p7_mult_21_n248, p7_mult_21_n247, p7_mult_21_n246, p7_mult_21_n245,
         p7_mult_21_n244, p7_mult_21_n243, p7_mult_21_n242, p7_mult_21_n241,
         p7_mult_21_n240, p7_mult_21_n239, p7_mult_21_n238, p7_mult_21_n237,
         p7_mult_21_n236, p7_mult_21_n235, p7_mult_21_n234, p7_mult_21_n233,
         p7_mult_21_n232, p7_mult_21_n231, p7_mult_21_n230, p7_mult_21_n229,
         p7_mult_21_n228, p7_mult_21_n227, p7_mult_21_n226, p7_mult_21_n225,
         p7_mult_21_n224, p7_mult_21_n223, p7_mult_21_n222, p7_mult_21_n221,
         p7_mult_21_n220, p7_mult_21_n219, p7_mult_21_n218, p7_mult_21_n217,
         p7_mult_21_n216, p7_mult_21_n215, p7_mult_21_n214, p7_mult_21_n213,
         p7_mult_21_n212, p7_mult_21_n211, p7_mult_21_n210, p7_mult_21_n209,
         p7_mult_21_n208, p7_mult_21_n207, p7_mult_21_n206, p7_mult_21_n205,
         p7_mult_21_n204, p7_mult_21_n203, p7_mult_21_n202, p7_mult_21_n201,
         p7_mult_21_n200, p7_mult_21_n199, p7_mult_21_n198, p7_mult_21_n197,
         p7_mult_21_n196, p7_mult_21_n195, p7_mult_21_n194, p7_mult_21_n193,
         p7_mult_21_n192, p7_mult_21_n191, p7_mult_21_n190, p7_mult_21_n189,
         p7_mult_21_n188, p7_mult_21_n187, p7_mult_21_n186, p7_mult_21_n185,
         p7_mult_21_n184, p7_mult_21_n183, p7_mult_21_n182, p7_mult_21_n181,
         p7_mult_21_n180, p7_mult_21_n179, p7_mult_21_n178, p7_mult_21_n177,
         p7_mult_21_n176, p7_mult_21_n175, p7_mult_21_n174, p7_mult_21_n173,
         p7_mult_21_n172, p7_mult_21_n171, p7_mult_21_n170, p7_mult_21_n169,
         p7_mult_21_n168, p7_mult_21_n167, p7_mult_21_n166, p7_mult_21_n165,
         p7_mult_21_n164, p7_mult_21_n163, p7_mult_21_n162, p7_mult_21_n149,
         p7_mult_21_n148, p7_mult_21_n147, p7_mult_21_n146, p7_mult_21_n145,
         p7_mult_21_n144, p7_mult_21_n143, p7_mult_21_n142, p7_mult_21_n141,
         p7_mult_21_n140, p7_mult_21_n139, p7_mult_21_n138, p7_mult_21_n137,
         p7_mult_21_n136, REG2_1_n89, REG2_1_n88, REG2_1_n87, REG2_1_n86,
         REG2_1_n85, REG2_1_n84, REG2_1_n83, REG2_1_n82, REG2_1_n81,
         REG2_1_n80, REG2_1_n79, REG2_1_n78, REG2_1_n77, REG2_1_n76,
         REG2_1_n75, REG2_1_n74, REG2_1_n73, REG2_1_n72, REG2_1_n71,
         REG2_1_n70, REG2_1_n69, REG2_1_n68, REG2_1_n67, REG2_1_n66,
         REG2_1_n65, REG2_1_n64, REG2_1_n63, REG2_1_n62, REG2_1_n61,
         REG2_1_n60, REG2_1_n59, REG2_1_n58, REG2_1_n57, REG2_1_n56,
         REG2_1_n55, REG2_1_n54, REG2_1_n53, REG2_1_n52, REG2_1_n51,
         REG2_1_n50, REG2_1_n49, REG2_1_n48, REG2_1_n47, REG2_1_n46,
         REG2_1_n45, REG2_1_n44, REG2_1_n43, REGISTER3_n89, REGISTER3_n88,
         REGISTER3_n87, REGISTER3_n86, REGISTER3_n85, REGISTER3_n84,
         REGISTER3_n83, REGISTER3_n82, REGISTER3_n81, REGISTER3_n80,
         REGISTER3_n79, REGISTER3_n78, REGISTER3_n77, REGISTER3_n76,
         REGISTER3_n75, REGISTER3_n74, REGISTER3_n73, REGISTER3_n72,
         REGISTER3_n71, REGISTER3_n70, REGISTER3_n69, REGISTER3_n68,
         REGISTER3_n67, REGISTER3_n66, REGISTER3_n65, REGISTER3_n64,
         REGISTER3_n63, REGISTER3_n62, REGISTER3_n61, REGISTER3_n60,
         REGISTER3_n59, REGISTER3_n58, REGISTER3_n57, REGISTER3_n56,
         REGISTER3_n55, REGISTER3_n54, REGISTER3_n53, REGISTER3_n52,
         REGISTER3_n51, REGISTER3_n50, REGISTER3_n49, REGISTER3_n48,
         REGISTER3_n47, REGISTER3_n46, REGISTER3_n45, REGISTER3_n44,
         REGISTER3_n43, p8_mult_21_n805, p8_mult_21_n804, p8_mult_21_n803,
         p8_mult_21_n802, p8_mult_21_n801, p8_mult_21_n800, p8_mult_21_n799,
         p8_mult_21_n798, p8_mult_21_n797, p8_mult_21_n796, p8_mult_21_n795,
         p8_mult_21_n794, p8_mult_21_n793, p8_mult_21_n792, p8_mult_21_n791,
         p8_mult_21_n790, p8_mult_21_n789, p8_mult_21_n788, p8_mult_21_n787,
         p8_mult_21_n786, p8_mult_21_n785, p8_mult_21_n784, p8_mult_21_n783,
         p8_mult_21_n782, p8_mult_21_n781, p8_mult_21_n780, p8_mult_21_n779,
         p8_mult_21_n778, p8_mult_21_n777, p8_mult_21_n776, p8_mult_21_n775,
         p8_mult_21_n774, p8_mult_21_n773, p8_mult_21_n772, p8_mult_21_n771,
         p8_mult_21_n770, p8_mult_21_n769, p8_mult_21_n768, p8_mult_21_n767,
         p8_mult_21_n766, p8_mult_21_n765, p8_mult_21_n764, p8_mult_21_n763,
         p8_mult_21_n762, p8_mult_21_n761, p8_mult_21_n760, p8_mult_21_n759,
         p8_mult_21_n758, p8_mult_21_n757, p8_mult_21_n756, p8_mult_21_n755,
         p8_mult_21_n754, p8_mult_21_n753, p8_mult_21_n752, p8_mult_21_n751,
         p8_mult_21_n750, p8_mult_21_n749, p8_mult_21_n748, p8_mult_21_n747,
         p8_mult_21_n746, p8_mult_21_n745, p8_mult_21_n744, p8_mult_21_n743,
         p8_mult_21_n742, p8_mult_21_n741, p8_mult_21_n740, p8_mult_21_n739,
         p8_mult_21_n738, p8_mult_21_n737, p8_mult_21_n736, p8_mult_21_n735,
         p8_mult_21_n734, p8_mult_21_n733, p8_mult_21_n732, p8_mult_21_n731,
         p8_mult_21_n730, p8_mult_21_n729, p8_mult_21_n728, p8_mult_21_n727,
         p8_mult_21_n726, p8_mult_21_n725, p8_mult_21_n724, p8_mult_21_n723,
         p8_mult_21_n722, p8_mult_21_n721, p8_mult_21_n720, p8_mult_21_n719,
         p8_mult_21_n718, p8_mult_21_n717, p8_mult_21_n716, p8_mult_21_n715,
         p8_mult_21_n714, p8_mult_21_n713, p8_mult_21_n712, p8_mult_21_n711,
         p8_mult_21_n710, p8_mult_21_n709, p8_mult_21_n708, p8_mult_21_n707,
         p8_mult_21_n706, p8_mult_21_n705, p8_mult_21_n704, p8_mult_21_n703,
         p8_mult_21_n702, p8_mult_21_n701, p8_mult_21_n700, p8_mult_21_n699,
         p8_mult_21_n698, p8_mult_21_n697, p8_mult_21_n696, p8_mult_21_n695,
         p8_mult_21_n694, p8_mult_21_n693, p8_mult_21_n692, p8_mult_21_n691,
         p8_mult_21_n690, p8_mult_21_n689, p8_mult_21_n688, p8_mult_21_n687,
         p8_mult_21_n686, p8_mult_21_n685, p8_mult_21_n684, p8_mult_21_n683,
         p8_mult_21_n682, p8_mult_21_n681, p8_mult_21_n680, p8_mult_21_n679,
         p8_mult_21_n678, p8_mult_21_n677, p8_mult_21_n676, p8_mult_21_n675,
         p8_mult_21_n674, p8_mult_21_n673, p8_mult_21_n672, p8_mult_21_n671,
         p8_mult_21_n670, p8_mult_21_n669, p8_mult_21_n668, p8_mult_21_n667,
         p8_mult_21_n666, p8_mult_21_n665, p8_mult_21_n664, p8_mult_21_n663,
         p8_mult_21_n662, p8_mult_21_n661, p8_mult_21_n660, p8_mult_21_n659,
         p8_mult_21_n658, p8_mult_21_n657, p8_mult_21_n656, p8_mult_21_n655,
         p8_mult_21_n654, p8_mult_21_n653, p8_mult_21_n652, p8_mult_21_n651,
         p8_mult_21_n650, p8_mult_21_n649, p8_mult_21_n648, p8_mult_21_n647,
         p8_mult_21_n646, p8_mult_21_n645, p8_mult_21_n644, p8_mult_21_n643,
         p8_mult_21_n642, p8_mult_21_n641, p8_mult_21_n640, p8_mult_21_n639,
         p8_mult_21_n638, p8_mult_21_n637, p8_mult_21_n636, p8_mult_21_n635,
         p8_mult_21_n419, p8_mult_21_n418, p8_mult_21_n417, p8_mult_21_n416,
         p8_mult_21_n415, p8_mult_21_n414, p8_mult_21_n413, p8_mult_21_n412,
         p8_mult_21_n411, p8_mult_21_n410, p8_mult_21_n409, p8_mult_21_n408,
         p8_mult_21_n406, p8_mult_21_n405, p8_mult_21_n404, p8_mult_21_n403,
         p8_mult_21_n402, p8_mult_21_n401, p8_mult_21_n400, p8_mult_21_n399,
         p8_mult_21_n398, p8_mult_21_n397, p8_mult_21_n396, p8_mult_21_n395,
         p8_mult_21_n394, p8_mult_21_n393, p8_mult_21_n392, p8_mult_21_n391,
         p8_mult_21_n390, p8_mult_21_n389, p8_mult_21_n388, p8_mult_21_n387,
         p8_mult_21_n386, p8_mult_21_n385, p8_mult_21_n384, p8_mult_21_n382,
         p8_mult_21_n381, p8_mult_21_n380, p8_mult_21_n379, p8_mult_21_n378,
         p8_mult_21_n377, p8_mult_21_n376, p8_mult_21_n375, p8_mult_21_n374,
         p8_mult_21_n373, p8_mult_21_n372, p8_mult_21_n371, p8_mult_21_n370,
         p8_mult_21_n369, p8_mult_21_n368, p8_mult_21_n367, p8_mult_21_n366,
         p8_mult_21_n365, p8_mult_21_n364, p8_mult_21_n363, p8_mult_21_n362,
         p8_mult_21_n361, p8_mult_21_n360, p8_mult_21_n359, p8_mult_21_n358,
         p8_mult_21_n357, p8_mult_21_n356, p8_mult_21_n355, p8_mult_21_n354,
         p8_mult_21_n353, p8_mult_21_n352, p8_mult_21_n351, p8_mult_21_n350,
         p8_mult_21_n349, p8_mult_21_n348, p8_mult_21_n346, p8_mult_21_n345,
         p8_mult_21_n344, p8_mult_21_n343, p8_mult_21_n342, p8_mult_21_n341,
         p8_mult_21_n340, p8_mult_21_n339, p8_mult_21_n338, p8_mult_21_n337,
         p8_mult_21_n336, p8_mult_21_n335, p8_mult_21_n334, p8_mult_21_n333,
         p8_mult_21_n332, p8_mult_21_n331, p8_mult_21_n330, p8_mult_21_n329,
         p8_mult_21_n328, p8_mult_21_n327, p8_mult_21_n326, p8_mult_21_n325,
         p8_mult_21_n321, p8_mult_21_n320, p8_mult_21_n319, p8_mult_21_n318,
         p8_mult_21_n317, p8_mult_21_n316, p8_mult_21_n315, p8_mult_21_n314,
         p8_mult_21_n313, p8_mult_21_n312, p8_mult_21_n311, p8_mult_21_n310,
         p8_mult_21_n309, p8_mult_21_n308, p8_mult_21_n307, p8_mult_21_n306,
         p8_mult_21_n305, p8_mult_21_n304, p8_mult_21_n303, p8_mult_21_n302,
         p8_mult_21_n301, p8_mult_21_n300, p8_mult_21_n299, p8_mult_21_n298,
         p8_mult_21_n297, p8_mult_21_n296, p8_mult_21_n295, p8_mult_21_n294,
         p8_mult_21_n293, p8_mult_21_n292, p8_mult_21_n291, p8_mult_21_n290,
         p8_mult_21_n289, p8_mult_21_n288, p8_mult_21_n287, p8_mult_21_n286,
         p8_mult_21_n285, p8_mult_21_n284, p8_mult_21_n283, p8_mult_21_n282,
         p8_mult_21_n281, p8_mult_21_n280, p8_mult_21_n279, p8_mult_21_n278,
         p8_mult_21_n277, p8_mult_21_n276, p8_mult_21_n275, p8_mult_21_n274,
         p8_mult_21_n273, p8_mult_21_n272, p8_mult_21_n271, p8_mult_21_n270,
         p8_mult_21_n269, p8_mult_21_n268, p8_mult_21_n267, p8_mult_21_n266,
         p8_mult_21_n265, p8_mult_21_n264, p8_mult_21_n263, p8_mult_21_n262,
         p8_mult_21_n261, p8_mult_21_n260, p8_mult_21_n259, p8_mult_21_n258,
         p8_mult_21_n257, p8_mult_21_n256, p8_mult_21_n255, p8_mult_21_n254,
         p8_mult_21_n253, p8_mult_21_n252, p8_mult_21_n251, p8_mult_21_n250,
         p8_mult_21_n249, p8_mult_21_n248, p8_mult_21_n247, p8_mult_21_n246,
         p8_mult_21_n245, p8_mult_21_n244, p8_mult_21_n243, p8_mult_21_n242,
         p8_mult_21_n241, p8_mult_21_n240, p8_mult_21_n239, p8_mult_21_n238,
         p8_mult_21_n237, p8_mult_21_n236, p8_mult_21_n235, p8_mult_21_n234,
         p8_mult_21_n233, p8_mult_21_n232, p8_mult_21_n231, p8_mult_21_n230,
         p8_mult_21_n229, p8_mult_21_n228, p8_mult_21_n227, p8_mult_21_n226,
         p8_mult_21_n225, p8_mult_21_n224, p8_mult_21_n223, p8_mult_21_n222,
         p8_mult_21_n221, p8_mult_21_n220, p8_mult_21_n219, p8_mult_21_n218,
         p8_mult_21_n217, p8_mult_21_n216, p8_mult_21_n215, p8_mult_21_n214,
         p8_mult_21_n213, p8_mult_21_n212, p8_mult_21_n211, p8_mult_21_n210,
         p8_mult_21_n209, p8_mult_21_n208, p8_mult_21_n207, p8_mult_21_n206,
         p8_mult_21_n205, p8_mult_21_n204, p8_mult_21_n203, p8_mult_21_n202,
         p8_mult_21_n201, p8_mult_21_n200, p8_mult_21_n199, p8_mult_21_n198,
         p8_mult_21_n197, p8_mult_21_n196, p8_mult_21_n195, p8_mult_21_n194,
         p8_mult_21_n193, p8_mult_21_n192, p8_mult_21_n191, p8_mult_21_n190,
         p8_mult_21_n189, p8_mult_21_n188, p8_mult_21_n187, p8_mult_21_n186,
         p8_mult_21_n185, p8_mult_21_n184, p8_mult_21_n183, p8_mult_21_n182,
         p8_mult_21_n181, p8_mult_21_n180, p8_mult_21_n179, p8_mult_21_n178,
         p8_mult_21_n177, p8_mult_21_n176, p8_mult_21_n175, p8_mult_21_n174,
         p8_mult_21_n173, p8_mult_21_n172, p8_mult_21_n171, p8_mult_21_n170,
         p8_mult_21_n169, p8_mult_21_n168, p8_mult_21_n167, p8_mult_21_n166,
         p8_mult_21_n165, p8_mult_21_n164, p8_mult_21_n163, p8_mult_21_n162,
         p8_mult_21_n149, p8_mult_21_n148, p8_mult_21_n147, p8_mult_21_n146,
         p8_mult_21_n145, p8_mult_21_n144, p8_mult_21_n143, p8_mult_21_n142,
         p8_mult_21_n141, p8_mult_21_n140, p8_mult_21_n139, p8_mult_21_n138,
         p8_mult_21_n137, p8_mult_21_n136, REG3_1_n89, REG3_1_n88, REG3_1_n87,
         REG3_1_n86, REG3_1_n85, REG3_1_n84, REG3_1_n83, REG3_1_n82,
         REG3_1_n81, REG3_1_n80, REG3_1_n79, REG3_1_n78, REG3_1_n77,
         REG3_1_n76, REG3_1_n75, REG3_1_n74, REG3_1_n73, REG3_1_n72,
         REG3_1_n71, REG3_1_n70, REG3_1_n69, REG3_1_n68, REG3_1_n67,
         REG3_1_n66, REG3_1_n65, REG3_1_n64, REG3_1_n63, REG3_1_n62,
         REG3_1_n61, REG3_1_n60, REG3_1_n59, REG3_1_n58, REG3_1_n57,
         REG3_1_n56, REG3_1_n55, REG3_1_n54, REG3_1_n53, REG3_1_n52,
         REG3_1_n51, REG3_1_n50, REG3_1_n49, REG3_1_n48, REG3_1_n47,
         REG3_1_n46, REG3_1_n45, REG3_1_n44, REG3_1_n43, REGISTER4_n89,
         REGISTER4_n88, REGISTER4_n87, REGISTER4_n86, REGISTER4_n85,
         REGISTER4_n84, REGISTER4_n83, REGISTER4_n82, REGISTER4_n81,
         REGISTER4_n80, REGISTER4_n79, REGISTER4_n78, REGISTER4_n77,
         REGISTER4_n76, REGISTER4_n75, REGISTER4_n74, REGISTER4_n73,
         REGISTER4_n72, REGISTER4_n71, REGISTER4_n70, REGISTER4_n69,
         REGISTER4_n68, REGISTER4_n67, REGISTER4_n66, REGISTER4_n65,
         REGISTER4_n64, REGISTER4_n63, REGISTER4_n62, REGISTER4_n61,
         REGISTER4_n60, REGISTER4_n59, REGISTER4_n58, REGISTER4_n57,
         REGISTER4_n56, REGISTER4_n55, REGISTER4_n54, REGISTER4_n53,
         REGISTER4_n52, REGISTER4_n51, REGISTER4_n50, REGISTER4_n49,
         REGISTER4_n48, REGISTER4_n47, REGISTER4_n46, REGISTER4_n45,
         REGISTER4_n44, REGISTER4_n43, p9_mult_21_n805, p9_mult_21_n804,
         p9_mult_21_n803, p9_mult_21_n802, p9_mult_21_n801, p9_mult_21_n800,
         p9_mult_21_n799, p9_mult_21_n798, p9_mult_21_n797, p9_mult_21_n796,
         p9_mult_21_n795, p9_mult_21_n794, p9_mult_21_n793, p9_mult_21_n792,
         p9_mult_21_n791, p9_mult_21_n790, p9_mult_21_n789, p9_mult_21_n788,
         p9_mult_21_n787, p9_mult_21_n786, p9_mult_21_n785, p9_mult_21_n784,
         p9_mult_21_n783, p9_mult_21_n782, p9_mult_21_n781, p9_mult_21_n780,
         p9_mult_21_n779, p9_mult_21_n778, p9_mult_21_n777, p9_mult_21_n776,
         p9_mult_21_n775, p9_mult_21_n774, p9_mult_21_n773, p9_mult_21_n772,
         p9_mult_21_n771, p9_mult_21_n770, p9_mult_21_n769, p9_mult_21_n768,
         p9_mult_21_n767, p9_mult_21_n766, p9_mult_21_n765, p9_mult_21_n764,
         p9_mult_21_n763, p9_mult_21_n762, p9_mult_21_n761, p9_mult_21_n760,
         p9_mult_21_n759, p9_mult_21_n758, p9_mult_21_n757, p9_mult_21_n756,
         p9_mult_21_n755, p9_mult_21_n754, p9_mult_21_n753, p9_mult_21_n752,
         p9_mult_21_n751, p9_mult_21_n750, p9_mult_21_n749, p9_mult_21_n748,
         p9_mult_21_n747, p9_mult_21_n746, p9_mult_21_n745, p9_mult_21_n744,
         p9_mult_21_n743, p9_mult_21_n742, p9_mult_21_n741, p9_mult_21_n740,
         p9_mult_21_n739, p9_mult_21_n738, p9_mult_21_n737, p9_mult_21_n736,
         p9_mult_21_n735, p9_mult_21_n734, p9_mult_21_n733, p9_mult_21_n732,
         p9_mult_21_n731, p9_mult_21_n730, p9_mult_21_n729, p9_mult_21_n728,
         p9_mult_21_n727, p9_mult_21_n726, p9_mult_21_n725, p9_mult_21_n724,
         p9_mult_21_n723, p9_mult_21_n722, p9_mult_21_n721, p9_mult_21_n720,
         p9_mult_21_n719, p9_mult_21_n718, p9_mult_21_n717, p9_mult_21_n716,
         p9_mult_21_n715, p9_mult_21_n714, p9_mult_21_n713, p9_mult_21_n712,
         p9_mult_21_n711, p9_mult_21_n710, p9_mult_21_n709, p9_mult_21_n708,
         p9_mult_21_n707, p9_mult_21_n706, p9_mult_21_n705, p9_mult_21_n704,
         p9_mult_21_n703, p9_mult_21_n702, p9_mult_21_n701, p9_mult_21_n700,
         p9_mult_21_n699, p9_mult_21_n698, p9_mult_21_n697, p9_mult_21_n696,
         p9_mult_21_n695, p9_mult_21_n694, p9_mult_21_n693, p9_mult_21_n692,
         p9_mult_21_n691, p9_mult_21_n690, p9_mult_21_n689, p9_mult_21_n688,
         p9_mult_21_n687, p9_mult_21_n686, p9_mult_21_n685, p9_mult_21_n684,
         p9_mult_21_n683, p9_mult_21_n682, p9_mult_21_n681, p9_mult_21_n680,
         p9_mult_21_n679, p9_mult_21_n678, p9_mult_21_n677, p9_mult_21_n676,
         p9_mult_21_n675, p9_mult_21_n674, p9_mult_21_n673, p9_mult_21_n672,
         p9_mult_21_n671, p9_mult_21_n670, p9_mult_21_n669, p9_mult_21_n668,
         p9_mult_21_n667, p9_mult_21_n666, p9_mult_21_n665, p9_mult_21_n664,
         p9_mult_21_n663, p9_mult_21_n662, p9_mult_21_n661, p9_mult_21_n660,
         p9_mult_21_n659, p9_mult_21_n658, p9_mult_21_n657, p9_mult_21_n656,
         p9_mult_21_n655, p9_mult_21_n654, p9_mult_21_n653, p9_mult_21_n652,
         p9_mult_21_n651, p9_mult_21_n650, p9_mult_21_n649, p9_mult_21_n648,
         p9_mult_21_n647, p9_mult_21_n646, p9_mult_21_n645, p9_mult_21_n644,
         p9_mult_21_n643, p9_mult_21_n642, p9_mult_21_n641, p9_mult_21_n640,
         p9_mult_21_n639, p9_mult_21_n638, p9_mult_21_n637, p9_mult_21_n636,
         p9_mult_21_n635, p9_mult_21_n419, p9_mult_21_n418, p9_mult_21_n417,
         p9_mult_21_n416, p9_mult_21_n415, p9_mult_21_n414, p9_mult_21_n413,
         p9_mult_21_n412, p9_mult_21_n411, p9_mult_21_n410, p9_mult_21_n409,
         p9_mult_21_n408, p9_mult_21_n406, p9_mult_21_n405, p9_mult_21_n404,
         p9_mult_21_n403, p9_mult_21_n402, p9_mult_21_n401, p9_mult_21_n400,
         p9_mult_21_n399, p9_mult_21_n398, p9_mult_21_n397, p9_mult_21_n396,
         p9_mult_21_n395, p9_mult_21_n394, p9_mult_21_n393, p9_mult_21_n392,
         p9_mult_21_n391, p9_mult_21_n390, p9_mult_21_n389, p9_mult_21_n388,
         p9_mult_21_n387, p9_mult_21_n386, p9_mult_21_n385, p9_mult_21_n384,
         p9_mult_21_n382, p9_mult_21_n381, p9_mult_21_n380, p9_mult_21_n379,
         p9_mult_21_n378, p9_mult_21_n377, p9_mult_21_n376, p9_mult_21_n375,
         p9_mult_21_n374, p9_mult_21_n373, p9_mult_21_n372, p9_mult_21_n371,
         p9_mult_21_n370, p9_mult_21_n369, p9_mult_21_n368, p9_mult_21_n367,
         p9_mult_21_n366, p9_mult_21_n365, p9_mult_21_n364, p9_mult_21_n363,
         p9_mult_21_n362, p9_mult_21_n361, p9_mult_21_n360, p9_mult_21_n359,
         p9_mult_21_n358, p9_mult_21_n357, p9_mult_21_n356, p9_mult_21_n355,
         p9_mult_21_n354, p9_mult_21_n353, p9_mult_21_n352, p9_mult_21_n351,
         p9_mult_21_n350, p9_mult_21_n349, p9_mult_21_n348, p9_mult_21_n346,
         p9_mult_21_n345, p9_mult_21_n344, p9_mult_21_n343, p9_mult_21_n342,
         p9_mult_21_n341, p9_mult_21_n340, p9_mult_21_n339, p9_mult_21_n338,
         p9_mult_21_n337, p9_mult_21_n336, p9_mult_21_n335, p9_mult_21_n334,
         p9_mult_21_n333, p9_mult_21_n332, p9_mult_21_n331, p9_mult_21_n330,
         p9_mult_21_n329, p9_mult_21_n328, p9_mult_21_n327, p9_mult_21_n326,
         p9_mult_21_n325, p9_mult_21_n321, p9_mult_21_n320, p9_mult_21_n319,
         p9_mult_21_n318, p9_mult_21_n317, p9_mult_21_n316, p9_mult_21_n315,
         p9_mult_21_n314, p9_mult_21_n313, p9_mult_21_n312, p9_mult_21_n311,
         p9_mult_21_n310, p9_mult_21_n309, p9_mult_21_n308, p9_mult_21_n307,
         p9_mult_21_n306, p9_mult_21_n305, p9_mult_21_n304, p9_mult_21_n303,
         p9_mult_21_n302, p9_mult_21_n301, p9_mult_21_n300, p9_mult_21_n299,
         p9_mult_21_n298, p9_mult_21_n297, p9_mult_21_n296, p9_mult_21_n295,
         p9_mult_21_n294, p9_mult_21_n293, p9_mult_21_n292, p9_mult_21_n291,
         p9_mult_21_n290, p9_mult_21_n289, p9_mult_21_n288, p9_mult_21_n287,
         p9_mult_21_n286, p9_mult_21_n285, p9_mult_21_n284, p9_mult_21_n283,
         p9_mult_21_n282, p9_mult_21_n281, p9_mult_21_n280, p9_mult_21_n279,
         p9_mult_21_n278, p9_mult_21_n277, p9_mult_21_n276, p9_mult_21_n275,
         p9_mult_21_n274, p9_mult_21_n273, p9_mult_21_n272, p9_mult_21_n271,
         p9_mult_21_n270, p9_mult_21_n269, p9_mult_21_n268, p9_mult_21_n267,
         p9_mult_21_n266, p9_mult_21_n265, p9_mult_21_n264, p9_mult_21_n263,
         p9_mult_21_n262, p9_mult_21_n261, p9_mult_21_n260, p9_mult_21_n259,
         p9_mult_21_n258, p9_mult_21_n257, p9_mult_21_n256, p9_mult_21_n255,
         p9_mult_21_n254, p9_mult_21_n253, p9_mult_21_n252, p9_mult_21_n251,
         p9_mult_21_n250, p9_mult_21_n249, p9_mult_21_n248, p9_mult_21_n247,
         p9_mult_21_n246, p9_mult_21_n245, p9_mult_21_n244, p9_mult_21_n243,
         p9_mult_21_n242, p9_mult_21_n241, p9_mult_21_n240, p9_mult_21_n239,
         p9_mult_21_n238, p9_mult_21_n237, p9_mult_21_n236, p9_mult_21_n235,
         p9_mult_21_n234, p9_mult_21_n233, p9_mult_21_n232, p9_mult_21_n231,
         p9_mult_21_n230, p9_mult_21_n229, p9_mult_21_n228, p9_mult_21_n227,
         p9_mult_21_n226, p9_mult_21_n225, p9_mult_21_n224, p9_mult_21_n223,
         p9_mult_21_n222, p9_mult_21_n221, p9_mult_21_n220, p9_mult_21_n219,
         p9_mult_21_n218, p9_mult_21_n217, p9_mult_21_n216, p9_mult_21_n215,
         p9_mult_21_n214, p9_mult_21_n213, p9_mult_21_n212, p9_mult_21_n211,
         p9_mult_21_n210, p9_mult_21_n209, p9_mult_21_n208, p9_mult_21_n207,
         p9_mult_21_n206, p9_mult_21_n205, p9_mult_21_n204, p9_mult_21_n203,
         p9_mult_21_n202, p9_mult_21_n201, p9_mult_21_n200, p9_mult_21_n199,
         p9_mult_21_n198, p9_mult_21_n197, p9_mult_21_n196, p9_mult_21_n195,
         p9_mult_21_n194, p9_mult_21_n193, p9_mult_21_n192, p9_mult_21_n191,
         p9_mult_21_n190, p9_mult_21_n189, p9_mult_21_n188, p9_mult_21_n187,
         p9_mult_21_n186, p9_mult_21_n185, p9_mult_21_n184, p9_mult_21_n183,
         p9_mult_21_n182, p9_mult_21_n181, p9_mult_21_n180, p9_mult_21_n179,
         p9_mult_21_n178, p9_mult_21_n177, p9_mult_21_n176, p9_mult_21_n175,
         p9_mult_21_n174, p9_mult_21_n173, p9_mult_21_n172, p9_mult_21_n171,
         p9_mult_21_n170, p9_mult_21_n169, p9_mult_21_n168, p9_mult_21_n167,
         p9_mult_21_n166, p9_mult_21_n165, p9_mult_21_n164, p9_mult_21_n163,
         p9_mult_21_n162, p9_mult_21_n149, p9_mult_21_n148, p9_mult_21_n147,
         p9_mult_21_n146, p9_mult_21_n145, p9_mult_21_n144, p9_mult_21_n143,
         p9_mult_21_n142, p9_mult_21_n141, p9_mult_21_n140, p9_mult_21_n139,
         p9_mult_21_n138, p9_mult_21_n137, p9_mult_21_n136, REG4_1_n89,
         REG4_1_n88, REG4_1_n87, REG4_1_n86, REG4_1_n85, REG4_1_n84,
         REG4_1_n83, REG4_1_n82, REG4_1_n81, REG4_1_n80, REG4_1_n79,
         REG4_1_n78, REG4_1_n77, REG4_1_n76, REG4_1_n75, REG4_1_n74,
         REG4_1_n73, REG4_1_n72, REG4_1_n71, REG4_1_n70, REG4_1_n69,
         REG4_1_n68, REG4_1_n67, REG4_1_n66, REG4_1_n65, REG4_1_n64,
         REG4_1_n63, REG4_1_n62, REG4_1_n61, REG4_1_n60, REG4_1_n59,
         REG4_1_n58, REG4_1_n57, REG4_1_n56, REG4_1_n55, REG4_1_n54,
         REG4_1_n53, REG4_1_n52, REG4_1_n51, REG4_1_n50, REG4_1_n49,
         REG4_1_n48, REG4_1_n47, REG4_1_n46, REG4_1_n45, REG4_1_n44,
         REG4_1_n43, p11_mult_21_n805, p11_mult_21_n804, p11_mult_21_n803,
         p11_mult_21_n802, p11_mult_21_n801, p11_mult_21_n800,
         p11_mult_21_n799, p11_mult_21_n798, p11_mult_21_n797,
         p11_mult_21_n796, p11_mult_21_n795, p11_mult_21_n794,
         p11_mult_21_n793, p11_mult_21_n792, p11_mult_21_n791,
         p11_mult_21_n790, p11_mult_21_n789, p11_mult_21_n788,
         p11_mult_21_n787, p11_mult_21_n786, p11_mult_21_n785,
         p11_mult_21_n784, p11_mult_21_n783, p11_mult_21_n782,
         p11_mult_21_n781, p11_mult_21_n780, p11_mult_21_n779,
         p11_mult_21_n778, p11_mult_21_n777, p11_mult_21_n776,
         p11_mult_21_n775, p11_mult_21_n774, p11_mult_21_n773,
         p11_mult_21_n772, p11_mult_21_n771, p11_mult_21_n770,
         p11_mult_21_n769, p11_mult_21_n768, p11_mult_21_n767,
         p11_mult_21_n766, p11_mult_21_n765, p11_mult_21_n764,
         p11_mult_21_n763, p11_mult_21_n762, p11_mult_21_n761,
         p11_mult_21_n760, p11_mult_21_n759, p11_mult_21_n758,
         p11_mult_21_n757, p11_mult_21_n756, p11_mult_21_n755,
         p11_mult_21_n754, p11_mult_21_n753, p11_mult_21_n752,
         p11_mult_21_n751, p11_mult_21_n750, p11_mult_21_n749,
         p11_mult_21_n748, p11_mult_21_n747, p11_mult_21_n746,
         p11_mult_21_n745, p11_mult_21_n744, p11_mult_21_n743,
         p11_mult_21_n742, p11_mult_21_n741, p11_mult_21_n740,
         p11_mult_21_n739, p11_mult_21_n738, p11_mult_21_n737,
         p11_mult_21_n736, p11_mult_21_n735, p11_mult_21_n734,
         p11_mult_21_n733, p11_mult_21_n732, p11_mult_21_n731,
         p11_mult_21_n730, p11_mult_21_n729, p11_mult_21_n728,
         p11_mult_21_n727, p11_mult_21_n726, p11_mult_21_n725,
         p11_mult_21_n724, p11_mult_21_n723, p11_mult_21_n722,
         p11_mult_21_n721, p11_mult_21_n720, p11_mult_21_n719,
         p11_mult_21_n718, p11_mult_21_n717, p11_mult_21_n716,
         p11_mult_21_n715, p11_mult_21_n714, p11_mult_21_n713,
         p11_mult_21_n712, p11_mult_21_n711, p11_mult_21_n710,
         p11_mult_21_n709, p11_mult_21_n708, p11_mult_21_n707,
         p11_mult_21_n706, p11_mult_21_n705, p11_mult_21_n704,
         p11_mult_21_n703, p11_mult_21_n702, p11_mult_21_n701,
         p11_mult_21_n700, p11_mult_21_n699, p11_mult_21_n698,
         p11_mult_21_n697, p11_mult_21_n696, p11_mult_21_n695,
         p11_mult_21_n694, p11_mult_21_n693, p11_mult_21_n692,
         p11_mult_21_n691, p11_mult_21_n690, p11_mult_21_n689,
         p11_mult_21_n688, p11_mult_21_n687, p11_mult_21_n686,
         p11_mult_21_n685, p11_mult_21_n684, p11_mult_21_n683,
         p11_mult_21_n682, p11_mult_21_n681, p11_mult_21_n680,
         p11_mult_21_n679, p11_mult_21_n678, p11_mult_21_n677,
         p11_mult_21_n676, p11_mult_21_n675, p11_mult_21_n674,
         p11_mult_21_n673, p11_mult_21_n672, p11_mult_21_n671,
         p11_mult_21_n670, p11_mult_21_n669, p11_mult_21_n668,
         p11_mult_21_n667, p11_mult_21_n666, p11_mult_21_n665,
         p11_mult_21_n664, p11_mult_21_n663, p11_mult_21_n662,
         p11_mult_21_n661, p11_mult_21_n660, p11_mult_21_n659,
         p11_mult_21_n658, p11_mult_21_n657, p11_mult_21_n656,
         p11_mult_21_n655, p11_mult_21_n654, p11_mult_21_n653,
         p11_mult_21_n652, p11_mult_21_n651, p11_mult_21_n650,
         p11_mult_21_n649, p11_mult_21_n648, p11_mult_21_n647,
         p11_mult_21_n646, p11_mult_21_n645, p11_mult_21_n644,
         p11_mult_21_n643, p11_mult_21_n642, p11_mult_21_n641,
         p11_mult_21_n640, p11_mult_21_n639, p11_mult_21_n638,
         p11_mult_21_n637, p11_mult_21_n636, p11_mult_21_n635,
         p11_mult_21_n419, p11_mult_21_n418, p11_mult_21_n417,
         p11_mult_21_n416, p11_mult_21_n415, p11_mult_21_n414,
         p11_mult_21_n413, p11_mult_21_n412, p11_mult_21_n411,
         p11_mult_21_n410, p11_mult_21_n409, p11_mult_21_n408,
         p11_mult_21_n406, p11_mult_21_n405, p11_mult_21_n404,
         p11_mult_21_n403, p11_mult_21_n402, p11_mult_21_n401,
         p11_mult_21_n400, p11_mult_21_n399, p11_mult_21_n398,
         p11_mult_21_n397, p11_mult_21_n396, p11_mult_21_n395,
         p11_mult_21_n394, p11_mult_21_n393, p11_mult_21_n392,
         p11_mult_21_n391, p11_mult_21_n390, p11_mult_21_n389,
         p11_mult_21_n388, p11_mult_21_n387, p11_mult_21_n386,
         p11_mult_21_n385, p11_mult_21_n384, p11_mult_21_n382,
         p11_mult_21_n381, p11_mult_21_n380, p11_mult_21_n379,
         p11_mult_21_n378, p11_mult_21_n377, p11_mult_21_n376,
         p11_mult_21_n375, p11_mult_21_n374, p11_mult_21_n373,
         p11_mult_21_n372, p11_mult_21_n371, p11_mult_21_n370,
         p11_mult_21_n369, p11_mult_21_n368, p11_mult_21_n367,
         p11_mult_21_n366, p11_mult_21_n365, p11_mult_21_n364,
         p11_mult_21_n363, p11_mult_21_n362, p11_mult_21_n361,
         p11_mult_21_n360, p11_mult_21_n359, p11_mult_21_n358,
         p11_mult_21_n357, p11_mult_21_n356, p11_mult_21_n355,
         p11_mult_21_n354, p11_mult_21_n353, p11_mult_21_n352,
         p11_mult_21_n351, p11_mult_21_n350, p11_mult_21_n349,
         p11_mult_21_n348, p11_mult_21_n346, p11_mult_21_n345,
         p11_mult_21_n344, p11_mult_21_n343, p11_mult_21_n342,
         p11_mult_21_n341, p11_mult_21_n340, p11_mult_21_n339,
         p11_mult_21_n338, p11_mult_21_n337, p11_mult_21_n336,
         p11_mult_21_n335, p11_mult_21_n334, p11_mult_21_n333,
         p11_mult_21_n332, p11_mult_21_n331, p11_mult_21_n330,
         p11_mult_21_n329, p11_mult_21_n328, p11_mult_21_n327,
         p11_mult_21_n326, p11_mult_21_n325, p11_mult_21_n321,
         p11_mult_21_n320, p11_mult_21_n319, p11_mult_21_n318,
         p11_mult_21_n317, p11_mult_21_n316, p11_mult_21_n315,
         p11_mult_21_n314, p11_mult_21_n313, p11_mult_21_n312,
         p11_mult_21_n311, p11_mult_21_n310, p11_mult_21_n309,
         p11_mult_21_n308, p11_mult_21_n307, p11_mult_21_n306,
         p11_mult_21_n305, p11_mult_21_n304, p11_mult_21_n303,
         p11_mult_21_n302, p11_mult_21_n301, p11_mult_21_n300,
         p11_mult_21_n299, p11_mult_21_n298, p11_mult_21_n297,
         p11_mult_21_n296, p11_mult_21_n295, p11_mult_21_n294,
         p11_mult_21_n293, p11_mult_21_n292, p11_mult_21_n291,
         p11_mult_21_n290, p11_mult_21_n289, p11_mult_21_n288,
         p11_mult_21_n287, p11_mult_21_n286, p11_mult_21_n285,
         p11_mult_21_n284, p11_mult_21_n283, p11_mult_21_n282,
         p11_mult_21_n281, p11_mult_21_n280, p11_mult_21_n279,
         p11_mult_21_n278, p11_mult_21_n277, p11_mult_21_n276,
         p11_mult_21_n275, p11_mult_21_n274, p11_mult_21_n273,
         p11_mult_21_n272, p11_mult_21_n271, p11_mult_21_n270,
         p11_mult_21_n269, p11_mult_21_n268, p11_mult_21_n267,
         p11_mult_21_n266, p11_mult_21_n265, p11_mult_21_n264,
         p11_mult_21_n263, p11_mult_21_n262, p11_mult_21_n261,
         p11_mult_21_n260, p11_mult_21_n259, p11_mult_21_n258,
         p11_mult_21_n257, p11_mult_21_n256, p11_mult_21_n255,
         p11_mult_21_n254, p11_mult_21_n253, p11_mult_21_n252,
         p11_mult_21_n251, p11_mult_21_n250, p11_mult_21_n249,
         p11_mult_21_n248, p11_mult_21_n247, p11_mult_21_n246,
         p11_mult_21_n245, p11_mult_21_n244, p11_mult_21_n243,
         p11_mult_21_n242, p11_mult_21_n241, p11_mult_21_n240,
         p11_mult_21_n239, p11_mult_21_n238, p11_mult_21_n237,
         p11_mult_21_n236, p11_mult_21_n235, p11_mult_21_n234,
         p11_mult_21_n233, p11_mult_21_n232, p11_mult_21_n231,
         p11_mult_21_n230, p11_mult_21_n229, p11_mult_21_n228,
         p11_mult_21_n227, p11_mult_21_n226, p11_mult_21_n225,
         p11_mult_21_n224, p11_mult_21_n223, p11_mult_21_n222,
         p11_mult_21_n221, p11_mult_21_n220, p11_mult_21_n219,
         p11_mult_21_n218, p11_mult_21_n217, p11_mult_21_n216,
         p11_mult_21_n215, p11_mult_21_n214, p11_mult_21_n213,
         p11_mult_21_n212, p11_mult_21_n211, p11_mult_21_n210,
         p11_mult_21_n209, p11_mult_21_n208, p11_mult_21_n207,
         p11_mult_21_n206, p11_mult_21_n205, p11_mult_21_n204,
         p11_mult_21_n203, p11_mult_21_n202, p11_mult_21_n201,
         p11_mult_21_n200, p11_mult_21_n199, p11_mult_21_n198,
         p11_mult_21_n197, p11_mult_21_n196, p11_mult_21_n195,
         p11_mult_21_n194, p11_mult_21_n193, p11_mult_21_n192,
         p11_mult_21_n191, p11_mult_21_n190, p11_mult_21_n189,
         p11_mult_21_n188, p11_mult_21_n187, p11_mult_21_n186,
         p11_mult_21_n185, p11_mult_21_n184, p11_mult_21_n183,
         p11_mult_21_n182, p11_mult_21_n181, p11_mult_21_n180,
         p11_mult_21_n179, p11_mult_21_n178, p11_mult_21_n177,
         p11_mult_21_n176, p11_mult_21_n175, p11_mult_21_n174,
         p11_mult_21_n173, p11_mult_21_n172, p11_mult_21_n171,
         p11_mult_21_n170, p11_mult_21_n169, p11_mult_21_n168,
         p11_mult_21_n167, p11_mult_21_n166, p11_mult_21_n165,
         p11_mult_21_n164, p11_mult_21_n163, p11_mult_21_n162,
         p11_mult_21_n149, p11_mult_21_n148, p11_mult_21_n147,
         p11_mult_21_n146, p11_mult_21_n145, p11_mult_21_n144,
         p11_mult_21_n143, p11_mult_21_n142, p11_mult_21_n141,
         p11_mult_21_n140, p11_mult_21_n139, p11_mult_21_n138,
         p11_mult_21_n137, p11_mult_21_n136, p10_mult_21_n805,
         p10_mult_21_n804, p10_mult_21_n803, p10_mult_21_n802,
         p10_mult_21_n801, p10_mult_21_n800, p10_mult_21_n799,
         p10_mult_21_n798, p10_mult_21_n797, p10_mult_21_n796,
         p10_mult_21_n795, p10_mult_21_n794, p10_mult_21_n793,
         p10_mult_21_n792, p10_mult_21_n791, p10_mult_21_n790,
         p10_mult_21_n789, p10_mult_21_n788, p10_mult_21_n787,
         p10_mult_21_n786, p10_mult_21_n785, p10_mult_21_n784,
         p10_mult_21_n783, p10_mult_21_n782, p10_mult_21_n781,
         p10_mult_21_n780, p10_mult_21_n779, p10_mult_21_n778,
         p10_mult_21_n777, p10_mult_21_n776, p10_mult_21_n775,
         p10_mult_21_n774, p10_mult_21_n773, p10_mult_21_n772,
         p10_mult_21_n771, p10_mult_21_n770, p10_mult_21_n769,
         p10_mult_21_n768, p10_mult_21_n767, p10_mult_21_n766,
         p10_mult_21_n765, p10_mult_21_n764, p10_mult_21_n763,
         p10_mult_21_n762, p10_mult_21_n761, p10_mult_21_n760,
         p10_mult_21_n759, p10_mult_21_n758, p10_mult_21_n757,
         p10_mult_21_n756, p10_mult_21_n755, p10_mult_21_n754,
         p10_mult_21_n753, p10_mult_21_n752, p10_mult_21_n751,
         p10_mult_21_n750, p10_mult_21_n749, p10_mult_21_n748,
         p10_mult_21_n747, p10_mult_21_n746, p10_mult_21_n745,
         p10_mult_21_n744, p10_mult_21_n743, p10_mult_21_n742,
         p10_mult_21_n741, p10_mult_21_n740, p10_mult_21_n739,
         p10_mult_21_n738, p10_mult_21_n737, p10_mult_21_n736,
         p10_mult_21_n735, p10_mult_21_n734, p10_mult_21_n733,
         p10_mult_21_n732, p10_mult_21_n731, p10_mult_21_n730,
         p10_mult_21_n729, p10_mult_21_n728, p10_mult_21_n727,
         p10_mult_21_n726, p10_mult_21_n725, p10_mult_21_n724,
         p10_mult_21_n723, p10_mult_21_n722, p10_mult_21_n721,
         p10_mult_21_n720, p10_mult_21_n719, p10_mult_21_n718,
         p10_mult_21_n717, p10_mult_21_n716, p10_mult_21_n715,
         p10_mult_21_n714, p10_mult_21_n713, p10_mult_21_n712,
         p10_mult_21_n711, p10_mult_21_n710, p10_mult_21_n709,
         p10_mult_21_n708, p10_mult_21_n707, p10_mult_21_n706,
         p10_mult_21_n705, p10_mult_21_n704, p10_mult_21_n703,
         p10_mult_21_n702, p10_mult_21_n701, p10_mult_21_n700,
         p10_mult_21_n699, p10_mult_21_n698, p10_mult_21_n697,
         p10_mult_21_n696, p10_mult_21_n695, p10_mult_21_n694,
         p10_mult_21_n693, p10_mult_21_n692, p10_mult_21_n691,
         p10_mult_21_n690, p10_mult_21_n689, p10_mult_21_n688,
         p10_mult_21_n687, p10_mult_21_n686, p10_mult_21_n685,
         p10_mult_21_n684, p10_mult_21_n683, p10_mult_21_n682,
         p10_mult_21_n681, p10_mult_21_n680, p10_mult_21_n679,
         p10_mult_21_n678, p10_mult_21_n677, p10_mult_21_n676,
         p10_mult_21_n675, p10_mult_21_n674, p10_mult_21_n673,
         p10_mult_21_n672, p10_mult_21_n671, p10_mult_21_n670,
         p10_mult_21_n669, p10_mult_21_n668, p10_mult_21_n667,
         p10_mult_21_n666, p10_mult_21_n665, p10_mult_21_n664,
         p10_mult_21_n663, p10_mult_21_n662, p10_mult_21_n661,
         p10_mult_21_n660, p10_mult_21_n659, p10_mult_21_n658,
         p10_mult_21_n657, p10_mult_21_n656, p10_mult_21_n655,
         p10_mult_21_n654, p10_mult_21_n653, p10_mult_21_n652,
         p10_mult_21_n651, p10_mult_21_n650, p10_mult_21_n649,
         p10_mult_21_n648, p10_mult_21_n647, p10_mult_21_n646,
         p10_mult_21_n645, p10_mult_21_n644, p10_mult_21_n643,
         p10_mult_21_n642, p10_mult_21_n641, p10_mult_21_n640,
         p10_mult_21_n639, p10_mult_21_n638, p10_mult_21_n637,
         p10_mult_21_n636, p10_mult_21_n635, p10_mult_21_n419,
         p10_mult_21_n418, p10_mult_21_n417, p10_mult_21_n416,
         p10_mult_21_n415, p10_mult_21_n414, p10_mult_21_n413,
         p10_mult_21_n412, p10_mult_21_n411, p10_mult_21_n410,
         p10_mult_21_n409, p10_mult_21_n408, p10_mult_21_n406,
         p10_mult_21_n405, p10_mult_21_n404, p10_mult_21_n403,
         p10_mult_21_n402, p10_mult_21_n401, p10_mult_21_n400,
         p10_mult_21_n399, p10_mult_21_n398, p10_mult_21_n397,
         p10_mult_21_n396, p10_mult_21_n395, p10_mult_21_n394,
         p10_mult_21_n393, p10_mult_21_n392, p10_mult_21_n391,
         p10_mult_21_n390, p10_mult_21_n389, p10_mult_21_n388,
         p10_mult_21_n387, p10_mult_21_n386, p10_mult_21_n385,
         p10_mult_21_n384, p10_mult_21_n382, p10_mult_21_n381,
         p10_mult_21_n380, p10_mult_21_n379, p10_mult_21_n378,
         p10_mult_21_n377, p10_mult_21_n376, p10_mult_21_n375,
         p10_mult_21_n374, p10_mult_21_n373, p10_mult_21_n372,
         p10_mult_21_n371, p10_mult_21_n370, p10_mult_21_n369,
         p10_mult_21_n368, p10_mult_21_n367, p10_mult_21_n366,
         p10_mult_21_n365, p10_mult_21_n364, p10_mult_21_n363,
         p10_mult_21_n362, p10_mult_21_n361, p10_mult_21_n360,
         p10_mult_21_n359, p10_mult_21_n358, p10_mult_21_n357,
         p10_mult_21_n356, p10_mult_21_n355, p10_mult_21_n354,
         p10_mult_21_n353, p10_mult_21_n352, p10_mult_21_n351,
         p10_mult_21_n350, p10_mult_21_n349, p10_mult_21_n348,
         p10_mult_21_n346, p10_mult_21_n345, p10_mult_21_n344,
         p10_mult_21_n343, p10_mult_21_n342, p10_mult_21_n341,
         p10_mult_21_n340, p10_mult_21_n339, p10_mult_21_n338,
         p10_mult_21_n337, p10_mult_21_n336, p10_mult_21_n335,
         p10_mult_21_n334, p10_mult_21_n333, p10_mult_21_n332,
         p10_mult_21_n331, p10_mult_21_n330, p10_mult_21_n329,
         p10_mult_21_n328, p10_mult_21_n327, p10_mult_21_n326,
         p10_mult_21_n325, p10_mult_21_n321, p10_mult_21_n320,
         p10_mult_21_n319, p10_mult_21_n318, p10_mult_21_n317,
         p10_mult_21_n316, p10_mult_21_n315, p10_mult_21_n314,
         p10_mult_21_n313, p10_mult_21_n312, p10_mult_21_n311,
         p10_mult_21_n310, p10_mult_21_n309, p10_mult_21_n308,
         p10_mult_21_n307, p10_mult_21_n306, p10_mult_21_n305,
         p10_mult_21_n304, p10_mult_21_n303, p10_mult_21_n302,
         p10_mult_21_n301, p10_mult_21_n300, p10_mult_21_n299,
         p10_mult_21_n298, p10_mult_21_n297, p10_mult_21_n296,
         p10_mult_21_n295, p10_mult_21_n294, p10_mult_21_n293,
         p10_mult_21_n292, p10_mult_21_n291, p10_mult_21_n290,
         p10_mult_21_n289, p10_mult_21_n288, p10_mult_21_n287,
         p10_mult_21_n286, p10_mult_21_n285, p10_mult_21_n284,
         p10_mult_21_n283, p10_mult_21_n282, p10_mult_21_n281,
         p10_mult_21_n280, p10_mult_21_n279, p10_mult_21_n278,
         p10_mult_21_n277, p10_mult_21_n276, p10_mult_21_n275,
         p10_mult_21_n274, p10_mult_21_n273, p10_mult_21_n272,
         p10_mult_21_n271, p10_mult_21_n270, p10_mult_21_n269,
         p10_mult_21_n268, p10_mult_21_n267, p10_mult_21_n266,
         p10_mult_21_n265, p10_mult_21_n264, p10_mult_21_n263,
         p10_mult_21_n262, p10_mult_21_n261, p10_mult_21_n260,
         p10_mult_21_n259, p10_mult_21_n258, p10_mult_21_n257,
         p10_mult_21_n256, p10_mult_21_n255, p10_mult_21_n254,
         p10_mult_21_n253, p10_mult_21_n252, p10_mult_21_n251,
         p10_mult_21_n250, p10_mult_21_n249, p10_mult_21_n248,
         p10_mult_21_n247, p10_mult_21_n246, p10_mult_21_n245,
         p10_mult_21_n244, p10_mult_21_n243, p10_mult_21_n242,
         p10_mult_21_n241, p10_mult_21_n240, p10_mult_21_n239,
         p10_mult_21_n238, p10_mult_21_n237, p10_mult_21_n236,
         p10_mult_21_n235, p10_mult_21_n234, p10_mult_21_n233,
         p10_mult_21_n232, p10_mult_21_n231, p10_mult_21_n230,
         p10_mult_21_n229, p10_mult_21_n228, p10_mult_21_n227,
         p10_mult_21_n226, p10_mult_21_n225, p10_mult_21_n224,
         p10_mult_21_n223, p10_mult_21_n222, p10_mult_21_n221,
         p10_mult_21_n220, p10_mult_21_n219, p10_mult_21_n218,
         p10_mult_21_n217, p10_mult_21_n216, p10_mult_21_n215,
         p10_mult_21_n214, p10_mult_21_n213, p10_mult_21_n212,
         p10_mult_21_n211, p10_mult_21_n210, p10_mult_21_n209,
         p10_mult_21_n208, p10_mult_21_n207, p10_mult_21_n206,
         p10_mult_21_n205, p10_mult_21_n204, p10_mult_21_n203,
         p10_mult_21_n202, p10_mult_21_n201, p10_mult_21_n200,
         p10_mult_21_n199, p10_mult_21_n198, p10_mult_21_n197,
         p10_mult_21_n196, p10_mult_21_n195, p10_mult_21_n194,
         p10_mult_21_n193, p10_mult_21_n192, p10_mult_21_n191,
         p10_mult_21_n190, p10_mult_21_n189, p10_mult_21_n188,
         p10_mult_21_n187, p10_mult_21_n186, p10_mult_21_n185,
         p10_mult_21_n184, p10_mult_21_n183, p10_mult_21_n182,
         p10_mult_21_n181, p10_mult_21_n180, p10_mult_21_n179,
         p10_mult_21_n178, p10_mult_21_n177, p10_mult_21_n176,
         p10_mult_21_n175, p10_mult_21_n174, p10_mult_21_n173,
         p10_mult_21_n172, p10_mult_21_n171, p10_mult_21_n170,
         p10_mult_21_n169, p10_mult_21_n168, p10_mult_21_n167,
         p10_mult_21_n166, p10_mult_21_n165, p10_mult_21_n164,
         p10_mult_21_n163, p10_mult_21_n162, p10_mult_21_n149,
         p10_mult_21_n148, p10_mult_21_n147, p10_mult_21_n146,
         p10_mult_21_n145, p10_mult_21_n144, p10_mult_21_n143,
         p10_mult_21_n142, p10_mult_21_n141, p10_mult_21_n140,
         p10_mult_21_n139, p10_mult_21_n138, p10_mult_21_n137,
         p10_mult_21_n136, SUB1_sub_1_root_sub_0_root_sub_21_2_carry_13_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_12_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_11_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_10_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_9_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_8_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_7_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_6_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_5_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_4_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_3_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_2_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_carry_1_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_13_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_12_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_11_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_10_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_9_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_8_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_7_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_6_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_5_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_4_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_3_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_2_,
         SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_1_, SUB1_N1, SUB1_N10,
         SUB1_N11, SUB1_N12, SUB1_N13, SUB1_N2, SUB1_N3, SUB1_N4, SUB1_N5,
         SUB1_N6, SUB1_N7, SUB1_N8, SUB1_N9,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_1_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_2_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_3_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_4_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_5_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_6_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_7_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_8_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_9_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_10_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_13_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_, s6_add_21_carry_1_,
         s6_add_21_carry_2_, s6_add_21_carry_3_, s6_add_21_carry_4_,
         s6_add_21_carry_5_, s6_add_21_carry_6_, s6_add_21_carry_7_,
         s6_add_21_carry_8_, s6_add_21_carry_9_, s6_add_21_carry_10_,
         s6_add_21_carry_11_, s6_add_21_carry_12_, s6_add_21_carry_13_,
         s7_add_21_carry_1_, s7_add_21_carry_2_, s7_add_21_carry_3_,
         s7_add_21_carry_4_, s7_add_21_carry_5_, s7_add_21_carry_6_,
         s7_add_21_carry_7_, s7_add_21_carry_8_, s7_add_21_carry_9_,
         s7_add_21_carry_10_, s7_add_21_carry_11_, s7_add_21_carry_12_,
         s7_add_21_carry_13_, s8_add_21_carry_1_, s8_add_21_carry_2_,
         s8_add_21_carry_3_, s8_add_21_carry_4_, s8_add_21_carry_5_,
         s8_add_21_carry_6_, s8_add_21_carry_7_, s8_add_21_carry_8_,
         s8_add_21_carry_9_, s8_add_21_carry_10_, s8_add_21_carry_11_,
         s8_add_21_carry_12_, s8_add_21_carry_13_, s9_add_21_carry_1_,
         s9_add_21_carry_2_, s9_add_21_carry_3_, s9_add_21_carry_4_,
         s9_add_21_carry_5_, s9_add_21_carry_6_, s9_add_21_carry_7_,
         s9_add_21_carry_8_, s9_add_21_carry_9_, s9_add_21_carry_10_,
         s9_add_21_carry_11_, s9_add_21_carry_12_, s9_add_21_carry_13_,
         REG11_n89, REG11_n88, REG11_n87, REG11_n86, REG11_n85, REG11_n84,
         REG11_n83, REG11_n82, REG11_n81, REG11_n80, REG11_n79, REG11_n78,
         REG11_n77, REG11_n76, REG11_n75, REG11_n74, REG11_n73, REG11_n72,
         REG11_n71, REG11_n70, REG11_n69, REG11_n68, REG11_n67, REG11_n66,
         REG11_n65, REG11_n64, REG11_n63, REG11_n62, REG11_n61, REG11_n60,
         REG11_n59, REG11_n58, REG11_n57, REG11_n56, REG11_n55, REG11_n54,
         REG11_n53, REG11_n52, REG11_n51, REG11_n50, REG11_n49, REG11_n48,
         REG11_n47, REG11_n46, REG11_n45, REG11_n44, REG11_n43, REG21_n89,
         REG21_n88, REG21_n87, REG21_n86, REG21_n85, REG21_n84, REG21_n83,
         REG21_n82, REG21_n81, REG21_n80, REG21_n79, REG21_n78, REG21_n77,
         REG21_n76, REG21_n75, REG21_n74, REG21_n73, REG21_n72, REG21_n71,
         REG21_n70, REG21_n69, REG21_n68, REG21_n67, REG21_n66, REG21_n65,
         REG21_n64, REG21_n63, REG21_n62, REG21_n61, REG21_n60, REG21_n59,
         REG21_n58, REG21_n57, REG21_n56, REG21_n55, REG21_n54, REG21_n53,
         REG21_n52, REG21_n51, REG21_n50, REG21_n49, REG21_n48, REG21_n47,
         REG21_n46, REG21_n45, REG21_n44, REG21_n43, REG31_n89, REG31_n88,
         REG31_n87, REG31_n86, REG31_n85, REG31_n84, REG31_n83, REG31_n82,
         REG31_n81, REG31_n80, REG31_n79, REG31_n78, REG31_n77, REG31_n76,
         REG31_n75, REG31_n74, REG31_n73, REG31_n72, REG31_n71, REG31_n70,
         REG31_n69, REG31_n68, REG31_n67, REG31_n66, REG31_n65, REG31_n64,
         REG31_n63, REG31_n62, REG31_n61, REG31_n60, REG31_n59, REG31_n58,
         REG31_n57, REG31_n56, REG31_n55, REG31_n54, REG31_n53, REG31_n52,
         REG31_n51, REG31_n50, REG31_n49, REG31_n48, REG31_n47, REG31_n46,
         REG31_n45, REG31_n44, REG31_n43, REG41_n89, REG41_n88, REG41_n87,
         REG41_n86, REG41_n85, REG41_n84, REG41_n83, REG41_n82, REG41_n81,
         REG41_n80, REG41_n79, REG41_n78, REG41_n77, REG41_n76, REG41_n75,
         REG41_n74, REG41_n73, REG41_n72, REG41_n71, REG41_n70, REG41_n69,
         REG41_n68, REG41_n67, REG41_n66, REG41_n65, REG41_n64, REG41_n63,
         REG41_n62, REG41_n61, REG41_n60, REG41_n59, REG41_n58, REG41_n57,
         REG41_n56, REG41_n55, REG41_n54, REG41_n53, REG41_n52, REG41_n51,
         REG41_n50, REG41_n49, REG41_n48, REG41_n47, REG41_n46, REG41_n45,
         REG41_n44, REG41_n43, REG51_n89, REG51_n88, REG51_n87, REG51_n86,
         REG51_n85, REG51_n84, REG51_n83, REG51_n82, REG51_n81, REG51_n80,
         REG51_n79, REG51_n78, REG51_n77, REG51_n76, REG51_n75, REG51_n74,
         REG51_n73, REG51_n72, REG51_n71, REG51_n70, REG51_n69, REG51_n68,
         REG51_n67, REG51_n66, REG51_n65, REG51_n64, REG51_n63, REG51_n62,
         REG51_n61, REG51_n60, REG51_n59, REG51_n58, REG51_n57, REG51_n56,
         REG51_n55, REG51_n54, REG51_n53, REG51_n52, REG51_n51, REG51_n50,
         REG51_n49, REG51_n48, REG51_n47, REG51_n46, REG51_n45, REG51_n44,
         REG51_n43, REG61_n89, REG61_n88, REG61_n87, REG61_n86, REG61_n85,
         REG61_n84, REG61_n83, REG61_n82, REG61_n81, REG61_n80, REG61_n79,
         REG61_n78, REG61_n77, REG61_n76, REG61_n75, REG61_n74, REG61_n73,
         REG61_n72, REG61_n71, REG61_n70, REG61_n69, REG61_n68, REG61_n67,
         REG61_n66, REG61_n65, REG61_n64, REG61_n63, REG61_n62, REG61_n61,
         REG61_n60, REG61_n59, REG61_n58, REG61_n57, REG61_n56, REG61_n55,
         REG61_n54, REG61_n53, REG61_n52, REG61_n51, REG61_n50, REG61_n49,
         REG61_n48, REG61_n47, REG61_n46, REG61_n45, REG61_n44, REG61_n43;
  wire   [13:0] w;
  wire   [13:0] reg1_reg;
  wire   [13:0] temp1;
  wire   [13:0] mul1_reg;
  wire   [13:0] reg2;
  wire   [13:0] reg2_reg;
  wire   [13:0] temp2;
  wire   [13:0] mul2_reg;
  wire   [13:0] reg3;
  wire   [13:0] reg3_reg;
  wire   [13:0] temp3;
  wire   [13:0] mul3_reg;
  wire   [13:0] reg5;
  wire   [13:0] reg4_reg;
  wire   [13:0] temp4;
  wire   [13:0] mul4_reg;
  wire   [13:0] temp6;
  wire   [13:0] reg4;
  wire   [13:0] temp5;
  wire   [13:0] reg6;
  wire   [13:0] reg7;
  wire   [13:0] fb;
  wire   [13:0] sig_ff1;
  wire   [13:0] sig_ff2;
  wire   [13:0] xin;

  DFFR_X1 xin_reg_13_ ( .D(n45), .CK(CLK), .RN(n48), .Q(xin[13]), .QN(n16) );
  DFFR_X1 xin_reg_12_ ( .D(n44), .CK(CLK), .RN(n48), .Q(xin[12]), .QN(n17) );
  DFFR_X1 xin_reg_11_ ( .D(n43), .CK(CLK), .RN(n48), .Q(xin[11]), .QN(n18) );
  DFFR_X1 xin_reg_10_ ( .D(n42), .CK(CLK), .RN(n48), .Q(xin[10]), .QN(n19) );
  DFFR_X1 xin_reg_9_ ( .D(n41), .CK(CLK), .RN(n48), .Q(xin[9]), .QN(n20) );
  DFFR_X1 xin_reg_8_ ( .D(n40), .CK(CLK), .RN(n48), .Q(xin[8]), .QN(n21) );
  DFFR_X1 xin_reg_7_ ( .D(n39), .CK(CLK), .RN(n48), .Q(xin[7]), .QN(n22) );
  DFFR_X1 xin_reg_6_ ( .D(n38), .CK(CLK), .RN(n48), .Q(xin[6]), .QN(n23) );
  DFFR_X1 xin_reg_5_ ( .D(n37), .CK(CLK), .RN(n48), .Q(xin[5]), .QN(n24) );
  DFFR_X1 xin_reg_4_ ( .D(n36), .CK(CLK), .RN(n48), .Q(xin[4]), .QN(n25) );
  DFFR_X1 xin_reg_3_ ( .D(n35), .CK(CLK), .RN(n48), .Q(xin[3]), .QN(n26) );
  DFFR_X1 xin_reg_2_ ( .D(n34), .CK(CLK), .RN(n48), .Q(xin[2]), .QN(n27) );
  DFFR_X1 xin_reg_1_ ( .D(n33), .CK(CLK), .RN(n48), .Q(xin[1]), .QN(n28) );
  DFFR_X1 xin_reg_0_ ( .D(n32), .CK(CLK), .RN(n48), .Q(xin[0]), .QN(n29) );
  DFFR_X1 VOUT_reg ( .D(n31), .CK(CLK), .RN(n48), .Q(VOUT), .QN(n30) );
  INV_X1 U33 ( .A(VIN), .ZN(n46) );
  OAI21_X1 U34 ( .B1(VIN), .B2(n29), .A(n2), .ZN(n32) );
  NAND2_X1 U35 ( .A1(VIN), .A2(DIN[0]), .ZN(n2) );
  OAI21_X1 U36 ( .B1(VIN), .B2(n27), .A(n4), .ZN(n34) );
  NAND2_X1 U37 ( .A1(DIN[2]), .A2(VIN), .ZN(n4) );
  OAI21_X1 U38 ( .B1(VIN), .B2(n26), .A(n5), .ZN(n35) );
  NAND2_X1 U39 ( .A1(DIN[3]), .A2(VIN), .ZN(n5) );
  OAI21_X1 U40 ( .B1(VIN), .B2(n28), .A(n3), .ZN(n33) );
  NAND2_X1 U41 ( .A1(DIN[1]), .A2(VIN), .ZN(n3) );
  OAI21_X1 U42 ( .B1(VIN), .B2(n25), .A(n6), .ZN(n36) );
  NAND2_X1 U43 ( .A1(DIN[4]), .A2(VIN), .ZN(n6) );
  OAI21_X1 U44 ( .B1(VIN), .B2(n24), .A(n7), .ZN(n37) );
  NAND2_X1 U45 ( .A1(DIN[5]), .A2(VIN), .ZN(n7) );
  OAI21_X1 U46 ( .B1(VIN), .B2(n23), .A(n8), .ZN(n38) );
  NAND2_X1 U47 ( .A1(DIN[6]), .A2(VIN), .ZN(n8) );
  OAI21_X1 U48 ( .B1(VIN), .B2(n22), .A(n9), .ZN(n39) );
  NAND2_X1 U49 ( .A1(DIN[7]), .A2(VIN), .ZN(n9) );
  OAI21_X1 U50 ( .B1(VIN), .B2(n21), .A(n10), .ZN(n40) );
  NAND2_X1 U51 ( .A1(DIN[8]), .A2(VIN), .ZN(n10) );
  OAI21_X1 U52 ( .B1(VIN), .B2(n20), .A(n11), .ZN(n41) );
  NAND2_X1 U53 ( .A1(DIN[9]), .A2(VIN), .ZN(n11) );
  OAI21_X1 U54 ( .B1(VIN), .B2(n19), .A(n12), .ZN(n42) );
  NAND2_X1 U55 ( .A1(DIN[10]), .A2(VIN), .ZN(n12) );
  OAI21_X1 U56 ( .B1(VIN), .B2(n18), .A(n13), .ZN(n43) );
  NAND2_X1 U57 ( .A1(DIN[11]), .A2(VIN), .ZN(n13) );
  OAI21_X1 U58 ( .B1(VIN), .B2(n17), .A(n14), .ZN(n44) );
  NAND2_X1 U59 ( .A1(DIN[12]), .A2(VIN), .ZN(n14) );
  OAI21_X1 U60 ( .B1(VIN), .B2(n16), .A(n15), .ZN(n45) );
  NAND2_X1 U61 ( .A1(DIN[13]), .A2(VIN), .ZN(n15) );
  NAND2_X1 U62 ( .A1(n30), .A2(n46), .ZN(n31) );
  BUF_X1 U63 ( .A(RST_n), .Z(n47) );
  BUF_X1 U64 ( .A(RST_n), .Z(n48) );
  NAND2_X1 REGISTER1_U34 ( .A1(w[13]), .A2(REGISTER1_n43), .ZN(REGISTER1_n14)
         );
  OAI21_X1 REGISTER1_U33 ( .B1(REGISTER1_n44), .B2(REGISTER1_n15), .A(
        REGISTER1_n14), .ZN(REGISTER1_n42) );
  NAND2_X1 REGISTER1_U32 ( .A1(w[6]), .A2(REGISTER1_n43), .ZN(REGISTER1_n7) );
  OAI21_X1 REGISTER1_U31 ( .B1(REGISTER1_n44), .B2(REGISTER1_n22), .A(
        REGISTER1_n7), .ZN(REGISTER1_n35) );
  NAND2_X1 REGISTER1_U30 ( .A1(w[5]), .A2(REGISTER1_n43), .ZN(REGISTER1_n6) );
  OAI21_X1 REGISTER1_U29 ( .B1(REGISTER1_n44), .B2(REGISTER1_n23), .A(
        REGISTER1_n6), .ZN(REGISTER1_n34) );
  NAND2_X1 REGISTER1_U28 ( .A1(w[4]), .A2(REGISTER1_n43), .ZN(REGISTER1_n5) );
  OAI21_X1 REGISTER1_U27 ( .B1(REGISTER1_n45), .B2(REGISTER1_n24), .A(
        REGISTER1_n5), .ZN(REGISTER1_n33) );
  NAND2_X1 REGISTER1_U26 ( .A1(w[3]), .A2(REGISTER1_n43), .ZN(REGISTER1_n4) );
  OAI21_X1 REGISTER1_U25 ( .B1(REGISTER1_n45), .B2(REGISTER1_n25), .A(
        REGISTER1_n4), .ZN(REGISTER1_n32) );
  NAND2_X1 REGISTER1_U24 ( .A1(w[2]), .A2(REGISTER1_n43), .ZN(REGISTER1_n3) );
  OAI21_X1 REGISTER1_U23 ( .B1(REGISTER1_n45), .B2(REGISTER1_n26), .A(
        REGISTER1_n3), .ZN(REGISTER1_n31) );
  NAND2_X1 REGISTER1_U22 ( .A1(w[1]), .A2(REGISTER1_n43), .ZN(REGISTER1_n2) );
  OAI21_X1 REGISTER1_U21 ( .B1(REGISTER1_n44), .B2(REGISTER1_n27), .A(
        REGISTER1_n2), .ZN(REGISTER1_n30) );
  NAND2_X1 REGISTER1_U20 ( .A1(w[8]), .A2(REGISTER1_n44), .ZN(REGISTER1_n9) );
  OAI21_X1 REGISTER1_U19 ( .B1(REGISTER1_n44), .B2(REGISTER1_n20), .A(
        REGISTER1_n9), .ZN(REGISTER1_n37) );
  NAND2_X1 REGISTER1_U18 ( .A1(w[12]), .A2(REGISTER1_n43), .ZN(REGISTER1_n13)
         );
  OAI21_X1 REGISTER1_U17 ( .B1(REGISTER1_n44), .B2(REGISTER1_n16), .A(
        REGISTER1_n13), .ZN(REGISTER1_n41) );
  NAND2_X1 REGISTER1_U16 ( .A1(w[11]), .A2(REGISTER1_n43), .ZN(REGISTER1_n12)
         );
  OAI21_X1 REGISTER1_U15 ( .B1(REGISTER1_n44), .B2(REGISTER1_n17), .A(
        REGISTER1_n12), .ZN(REGISTER1_n40) );
  NAND2_X1 REGISTER1_U14 ( .A1(w[10]), .A2(REGISTER1_n44), .ZN(REGISTER1_n11)
         );
  OAI21_X1 REGISTER1_U13 ( .B1(REGISTER1_n44), .B2(REGISTER1_n18), .A(
        REGISTER1_n11), .ZN(REGISTER1_n39) );
  NAND2_X1 REGISTER1_U12 ( .A1(w[9]), .A2(REGISTER1_n43), .ZN(REGISTER1_n10)
         );
  OAI21_X1 REGISTER1_U11 ( .B1(REGISTER1_n44), .B2(REGISTER1_n19), .A(
        REGISTER1_n10), .ZN(REGISTER1_n38) );
  NAND2_X1 REGISTER1_U10 ( .A1(w[7]), .A2(REGISTER1_n43), .ZN(REGISTER1_n8) );
  OAI21_X1 REGISTER1_U9 ( .B1(REGISTER1_n44), .B2(REGISTER1_n21), .A(
        REGISTER1_n8), .ZN(REGISTER1_n36) );
  NAND2_X1 REGISTER1_U8 ( .A1(w[0]), .A2(REGISTER1_n43), .ZN(REGISTER1_n1) );
  OAI21_X1 REGISTER1_U7 ( .B1(REGISTER1_n44), .B2(REGISTER1_n28), .A(
        REGISTER1_n1), .ZN(REGISTER1_n29) );
  BUF_X1 REGISTER1_U6 ( .A(n48), .Z(REGISTER1_n47) );
  BUF_X1 REGISTER1_U5 ( .A(n48), .Z(REGISTER1_n46) );
  BUF_X1 REGISTER1_U4 ( .A(VIN), .Z(REGISTER1_n45) );
  BUF_X1 REGISTER1_U3 ( .A(VIN), .Z(REGISTER1_n43) );
  BUF_X1 REGISTER1_U2 ( .A(VIN), .Z(REGISTER1_n44) );
  DFFR_X1 REGISTER1_q_reg_0_ ( .D(REGISTER1_n29), .CK(CLK), .RN(REGISTER1_n47), 
        .Q(reg1_reg[0]), .QN(REGISTER1_n28) );
  DFFR_X1 REGISTER1_q_reg_1_ ( .D(REGISTER1_n30), .CK(CLK), .RN(REGISTER1_n47), 
        .Q(reg1_reg[1]), .QN(REGISTER1_n27) );
  DFFR_X1 REGISTER1_q_reg_2_ ( .D(REGISTER1_n31), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[2]), .QN(REGISTER1_n26) );
  DFFR_X1 REGISTER1_q_reg_3_ ( .D(REGISTER1_n32), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[3]), .QN(REGISTER1_n25) );
  DFFR_X1 REGISTER1_q_reg_4_ ( .D(REGISTER1_n33), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[4]), .QN(REGISTER1_n24) );
  DFFR_X1 REGISTER1_q_reg_5_ ( .D(REGISTER1_n34), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[5]), .QN(REGISTER1_n23) );
  DFFR_X1 REGISTER1_q_reg_6_ ( .D(REGISTER1_n35), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[6]), .QN(REGISTER1_n22) );
  DFFR_X1 REGISTER1_q_reg_7_ ( .D(REGISTER1_n36), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[7]), .QN(REGISTER1_n21) );
  DFFR_X1 REGISTER1_q_reg_8_ ( .D(REGISTER1_n37), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[8]), .QN(REGISTER1_n20) );
  DFFR_X1 REGISTER1_q_reg_9_ ( .D(REGISTER1_n38), .CK(CLK), .RN(REGISTER1_n46), 
        .Q(reg1_reg[9]), .QN(REGISTER1_n19) );
  DFFR_X1 REGISTER1_q_reg_10_ ( .D(REGISTER1_n39), .CK(CLK), .RN(REGISTER1_n46), .Q(reg1_reg[10]), .QN(REGISTER1_n18) );
  DFFR_X1 REGISTER1_q_reg_11_ ( .D(REGISTER1_n40), .CK(CLK), .RN(REGISTER1_n46), .Q(reg1_reg[11]), .QN(REGISTER1_n17) );
  DFFR_X1 REGISTER1_q_reg_12_ ( .D(REGISTER1_n41), .CK(CLK), .RN(REGISTER1_n46), .Q(reg1_reg[12]), .QN(REGISTER1_n16) );
  DFFR_X1 REGISTER1_q_reg_13_ ( .D(REGISTER1_n42), .CK(CLK), .RN(REGISTER1_n46), .Q(reg1_reg[13]), .QN(REGISTER1_n15) );
  XOR2_X1 p6_mult_21_U691 ( .A(reg1_reg[2]), .B(reg1_reg[1]), .Z(
        p6_mult_21_n798) );
  INV_X1 p6_mult_21_U690 ( .A(reg1_reg[1]), .ZN(p6_mult_21_n655) );
  NOR2_X1 p6_mult_21_U689 ( .A1(p6_mult_21_n655), .A2(B0[1]), .ZN(
        p6_mult_21_n803) );
  INV_X1 p6_mult_21_U688 ( .A(p6_mult_21_n803), .ZN(p6_mult_21_n805) );
  NAND2_X1 p6_mult_21_U687 ( .A1(reg1_reg[1]), .A2(p6_mult_21_n643), .ZN(
        p6_mult_21_n641) );
  XNOR2_X1 p6_mult_21_U686 ( .A(B0[2]), .B(reg1_reg[1]), .ZN(p6_mult_21_n640)
         );
  OAI22_X1 p6_mult_21_U685 ( .A1(p6_mult_21_n805), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n640), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n804) );
  NAND2_X1 p6_mult_21_U684 ( .A1(p6_mult_21_n798), .A2(p6_mult_21_n804), .ZN(
        p6_mult_21_n801) );
  NAND2_X1 p6_mult_21_U683 ( .A1(p6_mult_21_n803), .A2(p6_mult_21_n804), .ZN(
        p6_mult_21_n802) );
  INV_X1 p6_mult_21_U682 ( .A(B0[0]), .ZN(p6_mult_21_n673) );
  MUX2_X1 p6_mult_21_U681 ( .A(p6_mult_21_n801), .B(p6_mult_21_n802), .S(
        p6_mult_21_n673), .Z(p6_mult_21_n800) );
  INV_X1 p6_mult_21_U680 ( .A(p6_mult_21_n800), .ZN(p6_mult_21_n795) );
  INV_X1 p6_mult_21_U679 ( .A(reg1_reg[3]), .ZN(p6_mult_21_n771) );
  XNOR2_X1 p6_mult_21_U678 ( .A(p6_mult_21_n771), .B(reg1_reg[2]), .ZN(
        p6_mult_21_n799) );
  NAND2_X1 p6_mult_21_U677 ( .A1(p6_mult_21_n658), .A2(p6_mult_21_n799), .ZN(
        p6_mult_21_n657) );
  NAND3_X1 p6_mult_21_U676 ( .A1(p6_mult_21_n798), .A2(p6_mult_21_n673), .A3(
        reg1_reg[3]), .ZN(p6_mult_21_n797) );
  OAI21_X1 p6_mult_21_U675 ( .B1(p6_mult_21_n771), .B2(p6_mult_21_n657), .A(
        p6_mult_21_n797), .ZN(p6_mult_21_n796) );
  AOI222_X1 p6_mult_21_U674 ( .A1(p6_mult_21_n795), .A2(p6_mult_21_n316), .B1(
        p6_mult_21_n796), .B2(p6_mult_21_n795), .C1(p6_mult_21_n796), .C2(
        p6_mult_21_n316), .ZN(p6_mult_21_n794) );
  INV_X1 p6_mult_21_U673 ( .A(p6_mult_21_n794), .ZN(p6_mult_21_n793) );
  AOI222_X1 p6_mult_21_U672 ( .A1(p6_mult_21_n793), .A2(p6_mult_21_n314), .B1(
        p6_mult_21_n793), .B2(p6_mult_21_n315), .C1(p6_mult_21_n315), .C2(
        p6_mult_21_n314), .ZN(p6_mult_21_n792) );
  INV_X1 p6_mult_21_U671 ( .A(p6_mult_21_n792), .ZN(p6_mult_21_n791) );
  AOI222_X1 p6_mult_21_U670 ( .A1(p6_mult_21_n791), .A2(p6_mult_21_n310), .B1(
        p6_mult_21_n791), .B2(p6_mult_21_n313), .C1(p6_mult_21_n313), .C2(
        p6_mult_21_n310), .ZN(p6_mult_21_n790) );
  INV_X1 p6_mult_21_U669 ( .A(p6_mult_21_n790), .ZN(p6_mult_21_n789) );
  AOI222_X1 p6_mult_21_U668 ( .A1(p6_mult_21_n789), .A2(p6_mult_21_n306), .B1(
        p6_mult_21_n789), .B2(p6_mult_21_n309), .C1(p6_mult_21_n309), .C2(
        p6_mult_21_n306), .ZN(p6_mult_21_n788) );
  INV_X1 p6_mult_21_U667 ( .A(p6_mult_21_n788), .ZN(p6_mult_21_n787) );
  AOI222_X1 p6_mult_21_U666 ( .A1(p6_mult_21_n787), .A2(p6_mult_21_n300), .B1(
        p6_mult_21_n787), .B2(p6_mult_21_n305), .C1(p6_mult_21_n305), .C2(
        p6_mult_21_n300), .ZN(p6_mult_21_n786) );
  INV_X1 p6_mult_21_U665 ( .A(p6_mult_21_n786), .ZN(p6_mult_21_n785) );
  AOI222_X1 p6_mult_21_U664 ( .A1(p6_mult_21_n785), .A2(p6_mult_21_n294), .B1(
        p6_mult_21_n785), .B2(p6_mult_21_n299), .C1(p6_mult_21_n299), .C2(
        p6_mult_21_n294), .ZN(p6_mult_21_n784) );
  INV_X1 p6_mult_21_U663 ( .A(p6_mult_21_n784), .ZN(p6_mult_21_n783) );
  AOI222_X1 p6_mult_21_U662 ( .A1(p6_mult_21_n783), .A2(p6_mult_21_n286), .B1(
        p6_mult_21_n783), .B2(p6_mult_21_n293), .C1(p6_mult_21_n293), .C2(
        p6_mult_21_n286), .ZN(p6_mult_21_n780) );
  INV_X1 p6_mult_21_U661 ( .A(p6_mult_21_n278), .ZN(p6_mult_21_n781) );
  INV_X1 p6_mult_21_U660 ( .A(p6_mult_21_n285), .ZN(p6_mult_21_n782) );
  OAI222_X1 p6_mult_21_U659 ( .A1(p6_mult_21_n780), .A2(p6_mult_21_n781), .B1(
        p6_mult_21_n780), .B2(p6_mult_21_n782), .C1(p6_mult_21_n782), .C2(
        p6_mult_21_n781), .ZN(p6_mult_21_n779) );
  AOI222_X1 p6_mult_21_U658 ( .A1(p6_mult_21_n779), .A2(p6_mult_21_n268), .B1(
        p6_mult_21_n779), .B2(p6_mult_21_n277), .C1(p6_mult_21_n277), .C2(
        p6_mult_21_n268), .ZN(p6_mult_21_n776) );
  INV_X1 p6_mult_21_U657 ( .A(p6_mult_21_n258), .ZN(p6_mult_21_n777) );
  INV_X1 p6_mult_21_U656 ( .A(p6_mult_21_n267), .ZN(p6_mult_21_n778) );
  OAI222_X1 p6_mult_21_U655 ( .A1(p6_mult_21_n776), .A2(p6_mult_21_n777), .B1(
        p6_mult_21_n776), .B2(p6_mult_21_n778), .C1(p6_mult_21_n778), .C2(
        p6_mult_21_n777), .ZN(p6_mult_21_n149) );
  XOR2_X1 p6_mult_21_U654 ( .A(B0[12]), .B(reg1_reg[13]), .Z(p6_mult_21_n757)
         );
  INV_X1 p6_mult_21_U653 ( .A(reg1_reg[11]), .ZN(p6_mult_21_n764) );
  INV_X1 p6_mult_21_U652 ( .A(reg1_reg[13]), .ZN(p6_mult_21_n766) );
  XNOR2_X1 p6_mult_21_U651 ( .A(p6_mult_21_n766), .B(reg1_reg[12]), .ZN(
        p6_mult_21_n775) );
  NAND2_X1 p6_mult_21_U650 ( .A1(p6_mult_21_n742), .A2(p6_mult_21_n775), .ZN(
        p6_mult_21_n744) );
  INV_X1 p6_mult_21_U649 ( .A(p6_mult_21_n744), .ZN(p6_mult_21_n637) );
  INV_X1 p6_mult_21_U648 ( .A(p6_mult_21_n742), .ZN(p6_mult_21_n638) );
  XNOR2_X1 p6_mult_21_U647 ( .A(B0[13]), .B(p6_mult_21_n766), .ZN(
        p6_mult_21_n639) );
  AOI22_X1 p6_mult_21_U646 ( .A1(p6_mult_21_n757), .A2(p6_mult_21_n637), .B1(
        p6_mult_21_n638), .B2(p6_mult_21_n639), .ZN(p6_mult_21_n162) );
  XNOR2_X1 p6_mult_21_U645 ( .A(B0[12]), .B(reg1_reg[11]), .ZN(p6_mult_21_n739) );
  INV_X1 p6_mult_21_U644 ( .A(reg1_reg[9]), .ZN(p6_mult_21_n762) );
  XNOR2_X1 p6_mult_21_U643 ( .A(p6_mult_21_n764), .B(reg1_reg[10]), .ZN(
        p6_mult_21_n774) );
  NAND2_X1 p6_mult_21_U642 ( .A1(p6_mult_21_n725), .A2(p6_mult_21_n774), .ZN(
        p6_mult_21_n727) );
  XNOR2_X1 p6_mult_21_U641 ( .A(B0[13]), .B(reg1_reg[11]), .ZN(p6_mult_21_n741) );
  OAI22_X1 p6_mult_21_U640 ( .A1(p6_mult_21_n739), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n741), .ZN(p6_mult_21_n167) );
  INV_X1 p6_mult_21_U639 ( .A(p6_mult_21_n167), .ZN(p6_mult_21_n168) );
  XNOR2_X1 p6_mult_21_U638 ( .A(B0[12]), .B(reg1_reg[9]), .ZN(p6_mult_21_n722)
         );
  INV_X1 p6_mult_21_U637 ( .A(reg1_reg[7]), .ZN(p6_mult_21_n760) );
  XNOR2_X1 p6_mult_21_U636 ( .A(p6_mult_21_n762), .B(reg1_reg[8]), .ZN(
        p6_mult_21_n773) );
  NAND2_X1 p6_mult_21_U635 ( .A1(p6_mult_21_n708), .A2(p6_mult_21_n773), .ZN(
        p6_mult_21_n710) );
  XNOR2_X1 p6_mult_21_U634 ( .A(B0[13]), .B(reg1_reg[9]), .ZN(p6_mult_21_n724)
         );
  OAI22_X1 p6_mult_21_U633 ( .A1(p6_mult_21_n722), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n724), .ZN(p6_mult_21_n177) );
  INV_X1 p6_mult_21_U632 ( .A(p6_mult_21_n177), .ZN(p6_mult_21_n178) );
  XNOR2_X1 p6_mult_21_U631 ( .A(B0[12]), .B(reg1_reg[7]), .ZN(p6_mult_21_n705)
         );
  INV_X1 p6_mult_21_U630 ( .A(reg1_reg[5]), .ZN(p6_mult_21_n758) );
  XNOR2_X1 p6_mult_21_U629 ( .A(p6_mult_21_n760), .B(reg1_reg[6]), .ZN(
        p6_mult_21_n772) );
  NAND2_X1 p6_mult_21_U628 ( .A1(p6_mult_21_n691), .A2(p6_mult_21_n772), .ZN(
        p6_mult_21_n693) );
  XNOR2_X1 p6_mult_21_U627 ( .A(B0[13]), .B(reg1_reg[7]), .ZN(p6_mult_21_n707)
         );
  OAI22_X1 p6_mult_21_U626 ( .A1(p6_mult_21_n705), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n707), .ZN(p6_mult_21_n191) );
  INV_X1 p6_mult_21_U625 ( .A(p6_mult_21_n191), .ZN(p6_mult_21_n192) );
  XNOR2_X1 p6_mult_21_U624 ( .A(B0[12]), .B(reg1_reg[5]), .ZN(p6_mult_21_n688)
         );
  XNOR2_X1 p6_mult_21_U623 ( .A(p6_mult_21_n758), .B(reg1_reg[4]), .ZN(
        p6_mult_21_n770) );
  NAND2_X1 p6_mult_21_U622 ( .A1(p6_mult_21_n674), .A2(p6_mult_21_n770), .ZN(
        p6_mult_21_n676) );
  XNOR2_X1 p6_mult_21_U621 ( .A(B0[13]), .B(reg1_reg[5]), .ZN(p6_mult_21_n690)
         );
  OAI22_X1 p6_mult_21_U620 ( .A1(p6_mult_21_n688), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n690), .ZN(p6_mult_21_n209) );
  INV_X1 p6_mult_21_U619 ( .A(p6_mult_21_n209), .ZN(p6_mult_21_n210) );
  XNOR2_X1 p6_mult_21_U618 ( .A(B0[12]), .B(reg1_reg[3]), .ZN(p6_mult_21_n670)
         );
  XNOR2_X1 p6_mult_21_U617 ( .A(B0[13]), .B(reg1_reg[3]), .ZN(p6_mult_21_n672)
         );
  OAI22_X1 p6_mult_21_U616 ( .A1(p6_mult_21_n670), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n672), .ZN(p6_mult_21_n231) );
  INV_X1 p6_mult_21_U615 ( .A(p6_mult_21_n231), .ZN(p6_mult_21_n232) );
  XNOR2_X1 p6_mult_21_U614 ( .A(B0[3]), .B(reg1_reg[11]), .ZN(p6_mult_21_n730)
         );
  XNOR2_X1 p6_mult_21_U613 ( .A(B0[4]), .B(reg1_reg[11]), .ZN(p6_mult_21_n731)
         );
  OAI22_X1 p6_mult_21_U612 ( .A1(p6_mult_21_n730), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n731), .ZN(p6_mult_21_n768) );
  XNOR2_X1 p6_mult_21_U611 ( .A(B0[9]), .B(reg1_reg[5]), .ZN(p6_mult_21_n685)
         );
  XNOR2_X1 p6_mult_21_U610 ( .A(B0[10]), .B(reg1_reg[5]), .ZN(p6_mult_21_n686)
         );
  OAI22_X1 p6_mult_21_U609 ( .A1(p6_mult_21_n685), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n686), .ZN(p6_mult_21_n769) );
  OR2_X1 p6_mult_21_U608 ( .A1(p6_mult_21_n768), .A2(p6_mult_21_n769), .ZN(
        p6_mult_21_n243) );
  XNOR2_X1 p6_mult_21_U607 ( .A(p6_mult_21_n768), .B(p6_mult_21_n769), .ZN(
        p6_mult_21_n244) );
  NAND3_X1 p6_mult_21_U606 ( .A1(p6_mult_21_n638), .A2(p6_mult_21_n673), .A3(
        reg1_reg[13]), .ZN(p6_mult_21_n767) );
  OAI21_X1 p6_mult_21_U605 ( .B1(p6_mult_21_n766), .B2(p6_mult_21_n744), .A(
        p6_mult_21_n767), .ZN(p6_mult_21_n317) );
  OR3_X1 p6_mult_21_U604 ( .A1(p6_mult_21_n725), .A2(B0[0]), .A3(
        p6_mult_21_n764), .ZN(p6_mult_21_n765) );
  OAI21_X1 p6_mult_21_U603 ( .B1(p6_mult_21_n764), .B2(p6_mult_21_n727), .A(
        p6_mult_21_n765), .ZN(p6_mult_21_n318) );
  OR3_X1 p6_mult_21_U602 ( .A1(p6_mult_21_n708), .A2(B0[0]), .A3(
        p6_mult_21_n762), .ZN(p6_mult_21_n763) );
  OAI21_X1 p6_mult_21_U601 ( .B1(p6_mult_21_n762), .B2(p6_mult_21_n710), .A(
        p6_mult_21_n763), .ZN(p6_mult_21_n319) );
  OR3_X1 p6_mult_21_U600 ( .A1(p6_mult_21_n691), .A2(B0[0]), .A3(
        p6_mult_21_n760), .ZN(p6_mult_21_n761) );
  OAI21_X1 p6_mult_21_U599 ( .B1(p6_mult_21_n760), .B2(p6_mult_21_n693), .A(
        p6_mult_21_n761), .ZN(p6_mult_21_n320) );
  OR3_X1 p6_mult_21_U598 ( .A1(p6_mult_21_n674), .A2(B0[0]), .A3(
        p6_mult_21_n758), .ZN(p6_mult_21_n759) );
  OAI21_X1 p6_mult_21_U597 ( .B1(p6_mult_21_n758), .B2(p6_mult_21_n676), .A(
        p6_mult_21_n759), .ZN(p6_mult_21_n321) );
  XNOR2_X1 p6_mult_21_U596 ( .A(B0[11]), .B(reg1_reg[13]), .ZN(p6_mult_21_n755) );
  INV_X1 p6_mult_21_U595 ( .A(p6_mult_21_n757), .ZN(p6_mult_21_n756) );
  OAI22_X1 p6_mult_21_U594 ( .A1(p6_mult_21_n755), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n756), .ZN(p6_mult_21_n325) );
  XNOR2_X1 p6_mult_21_U593 ( .A(B0[10]), .B(reg1_reg[13]), .ZN(p6_mult_21_n754) );
  OAI22_X1 p6_mult_21_U592 ( .A1(p6_mult_21_n754), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n755), .ZN(p6_mult_21_n326) );
  XNOR2_X1 p6_mult_21_U591 ( .A(B0[9]), .B(reg1_reg[13]), .ZN(p6_mult_21_n753)
         );
  OAI22_X1 p6_mult_21_U590 ( .A1(p6_mult_21_n753), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n754), .ZN(p6_mult_21_n327) );
  XNOR2_X1 p6_mult_21_U589 ( .A(B0[8]), .B(reg1_reg[13]), .ZN(p6_mult_21_n752)
         );
  OAI22_X1 p6_mult_21_U588 ( .A1(p6_mult_21_n752), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n753), .ZN(p6_mult_21_n328) );
  XNOR2_X1 p6_mult_21_U587 ( .A(B0[7]), .B(reg1_reg[13]), .ZN(p6_mult_21_n751)
         );
  OAI22_X1 p6_mult_21_U586 ( .A1(p6_mult_21_n751), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n752), .ZN(p6_mult_21_n329) );
  XNOR2_X1 p6_mult_21_U585 ( .A(B0[6]), .B(reg1_reg[13]), .ZN(p6_mult_21_n750)
         );
  OAI22_X1 p6_mult_21_U584 ( .A1(p6_mult_21_n750), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n751), .ZN(p6_mult_21_n330) );
  XNOR2_X1 p6_mult_21_U583 ( .A(B0[5]), .B(reg1_reg[13]), .ZN(p6_mult_21_n749)
         );
  OAI22_X1 p6_mult_21_U582 ( .A1(p6_mult_21_n749), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n750), .ZN(p6_mult_21_n331) );
  XNOR2_X1 p6_mult_21_U581 ( .A(B0[4]), .B(reg1_reg[13]), .ZN(p6_mult_21_n748)
         );
  OAI22_X1 p6_mult_21_U580 ( .A1(p6_mult_21_n748), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n749), .ZN(p6_mult_21_n332) );
  XNOR2_X1 p6_mult_21_U579 ( .A(B0[3]), .B(reg1_reg[13]), .ZN(p6_mult_21_n747)
         );
  OAI22_X1 p6_mult_21_U578 ( .A1(p6_mult_21_n747), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n748), .ZN(p6_mult_21_n333) );
  XNOR2_X1 p6_mult_21_U577 ( .A(B0[2]), .B(reg1_reg[13]), .ZN(p6_mult_21_n746)
         );
  OAI22_X1 p6_mult_21_U576 ( .A1(p6_mult_21_n746), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n747), .ZN(p6_mult_21_n334) );
  XNOR2_X1 p6_mult_21_U575 ( .A(B0[1]), .B(reg1_reg[13]), .ZN(p6_mult_21_n745)
         );
  OAI22_X1 p6_mult_21_U574 ( .A1(p6_mult_21_n745), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n746), .ZN(p6_mult_21_n335) );
  XNOR2_X1 p6_mult_21_U573 ( .A(reg1_reg[13]), .B(B0[0]), .ZN(p6_mult_21_n743)
         );
  OAI22_X1 p6_mult_21_U572 ( .A1(p6_mult_21_n743), .A2(p6_mult_21_n744), .B1(
        p6_mult_21_n742), .B2(p6_mult_21_n745), .ZN(p6_mult_21_n336) );
  NOR2_X1 p6_mult_21_U571 ( .A1(p6_mult_21_n673), .A2(p6_mult_21_n742), .ZN(
        p6_mult_21_n337) );
  AOI21_X1 p6_mult_21_U570 ( .B1(p6_mult_21_n727), .B2(p6_mult_21_n725), .A(
        p6_mult_21_n741), .ZN(p6_mult_21_n740) );
  INV_X1 p6_mult_21_U569 ( .A(p6_mult_21_n740), .ZN(p6_mult_21_n338) );
  XNOR2_X1 p6_mult_21_U568 ( .A(B0[11]), .B(reg1_reg[11]), .ZN(p6_mult_21_n738) );
  OAI22_X1 p6_mult_21_U567 ( .A1(p6_mult_21_n738), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n739), .ZN(p6_mult_21_n339) );
  XNOR2_X1 p6_mult_21_U566 ( .A(B0[10]), .B(reg1_reg[11]), .ZN(p6_mult_21_n737) );
  OAI22_X1 p6_mult_21_U565 ( .A1(p6_mult_21_n737), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n738), .ZN(p6_mult_21_n340) );
  XNOR2_X1 p6_mult_21_U564 ( .A(B0[9]), .B(reg1_reg[11]), .ZN(p6_mult_21_n736)
         );
  OAI22_X1 p6_mult_21_U563 ( .A1(p6_mult_21_n736), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n737), .ZN(p6_mult_21_n341) );
  XNOR2_X1 p6_mult_21_U562 ( .A(B0[8]), .B(reg1_reg[11]), .ZN(p6_mult_21_n735)
         );
  OAI22_X1 p6_mult_21_U561 ( .A1(p6_mult_21_n735), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n736), .ZN(p6_mult_21_n342) );
  XNOR2_X1 p6_mult_21_U560 ( .A(B0[7]), .B(reg1_reg[11]), .ZN(p6_mult_21_n734)
         );
  OAI22_X1 p6_mult_21_U559 ( .A1(p6_mult_21_n734), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n735), .ZN(p6_mult_21_n343) );
  XNOR2_X1 p6_mult_21_U558 ( .A(B0[6]), .B(reg1_reg[11]), .ZN(p6_mult_21_n733)
         );
  OAI22_X1 p6_mult_21_U557 ( .A1(p6_mult_21_n733), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n734), .ZN(p6_mult_21_n344) );
  XNOR2_X1 p6_mult_21_U556 ( .A(B0[5]), .B(reg1_reg[11]), .ZN(p6_mult_21_n732)
         );
  OAI22_X1 p6_mult_21_U555 ( .A1(p6_mult_21_n732), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n733), .ZN(p6_mult_21_n345) );
  OAI22_X1 p6_mult_21_U554 ( .A1(p6_mult_21_n731), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n732), .ZN(p6_mult_21_n346) );
  XNOR2_X1 p6_mult_21_U553 ( .A(B0[2]), .B(reg1_reg[11]), .ZN(p6_mult_21_n729)
         );
  OAI22_X1 p6_mult_21_U552 ( .A1(p6_mult_21_n729), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n730), .ZN(p6_mult_21_n348) );
  XNOR2_X1 p6_mult_21_U551 ( .A(B0[1]), .B(reg1_reg[11]), .ZN(p6_mult_21_n728)
         );
  OAI22_X1 p6_mult_21_U550 ( .A1(p6_mult_21_n728), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n729), .ZN(p6_mult_21_n349) );
  XNOR2_X1 p6_mult_21_U549 ( .A(reg1_reg[11]), .B(B0[0]), .ZN(p6_mult_21_n726)
         );
  OAI22_X1 p6_mult_21_U548 ( .A1(p6_mult_21_n726), .A2(p6_mult_21_n727), .B1(
        p6_mult_21_n725), .B2(p6_mult_21_n728), .ZN(p6_mult_21_n350) );
  NOR2_X1 p6_mult_21_U547 ( .A1(p6_mult_21_n673), .A2(p6_mult_21_n725), .ZN(
        p6_mult_21_n351) );
  AOI21_X1 p6_mult_21_U546 ( .B1(p6_mult_21_n710), .B2(p6_mult_21_n708), .A(
        p6_mult_21_n724), .ZN(p6_mult_21_n723) );
  INV_X1 p6_mult_21_U545 ( .A(p6_mult_21_n723), .ZN(p6_mult_21_n352) );
  XNOR2_X1 p6_mult_21_U544 ( .A(B0[11]), .B(reg1_reg[9]), .ZN(p6_mult_21_n721)
         );
  OAI22_X1 p6_mult_21_U543 ( .A1(p6_mult_21_n721), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n722), .ZN(p6_mult_21_n353) );
  XNOR2_X1 p6_mult_21_U542 ( .A(B0[10]), .B(reg1_reg[9]), .ZN(p6_mult_21_n720)
         );
  OAI22_X1 p6_mult_21_U541 ( .A1(p6_mult_21_n720), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n721), .ZN(p6_mult_21_n354) );
  XNOR2_X1 p6_mult_21_U540 ( .A(B0[9]), .B(reg1_reg[9]), .ZN(p6_mult_21_n719)
         );
  OAI22_X1 p6_mult_21_U539 ( .A1(p6_mult_21_n719), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n720), .ZN(p6_mult_21_n355) );
  XNOR2_X1 p6_mult_21_U538 ( .A(B0[8]), .B(reg1_reg[9]), .ZN(p6_mult_21_n718)
         );
  OAI22_X1 p6_mult_21_U537 ( .A1(p6_mult_21_n718), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n719), .ZN(p6_mult_21_n356) );
  XNOR2_X1 p6_mult_21_U536 ( .A(B0[7]), .B(reg1_reg[9]), .ZN(p6_mult_21_n717)
         );
  OAI22_X1 p6_mult_21_U535 ( .A1(p6_mult_21_n717), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n718), .ZN(p6_mult_21_n357) );
  XNOR2_X1 p6_mult_21_U534 ( .A(B0[6]), .B(reg1_reg[9]), .ZN(p6_mult_21_n716)
         );
  OAI22_X1 p6_mult_21_U533 ( .A1(p6_mult_21_n716), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n717), .ZN(p6_mult_21_n358) );
  XNOR2_X1 p6_mult_21_U532 ( .A(B0[5]), .B(reg1_reg[9]), .ZN(p6_mult_21_n715)
         );
  OAI22_X1 p6_mult_21_U531 ( .A1(p6_mult_21_n715), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n716), .ZN(p6_mult_21_n359) );
  XNOR2_X1 p6_mult_21_U530 ( .A(B0[4]), .B(reg1_reg[9]), .ZN(p6_mult_21_n714)
         );
  OAI22_X1 p6_mult_21_U529 ( .A1(p6_mult_21_n714), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n715), .ZN(p6_mult_21_n360) );
  XNOR2_X1 p6_mult_21_U528 ( .A(B0[3]), .B(reg1_reg[9]), .ZN(p6_mult_21_n713)
         );
  OAI22_X1 p6_mult_21_U527 ( .A1(p6_mult_21_n713), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n714), .ZN(p6_mult_21_n361) );
  XNOR2_X1 p6_mult_21_U526 ( .A(B0[2]), .B(reg1_reg[9]), .ZN(p6_mult_21_n712)
         );
  OAI22_X1 p6_mult_21_U525 ( .A1(p6_mult_21_n712), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n713), .ZN(p6_mult_21_n362) );
  XNOR2_X1 p6_mult_21_U524 ( .A(B0[1]), .B(reg1_reg[9]), .ZN(p6_mult_21_n711)
         );
  OAI22_X1 p6_mult_21_U523 ( .A1(p6_mult_21_n711), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n712), .ZN(p6_mult_21_n363) );
  XNOR2_X1 p6_mult_21_U522 ( .A(reg1_reg[9]), .B(B0[0]), .ZN(p6_mult_21_n709)
         );
  OAI22_X1 p6_mult_21_U521 ( .A1(p6_mult_21_n709), .A2(p6_mult_21_n710), .B1(
        p6_mult_21_n708), .B2(p6_mult_21_n711), .ZN(p6_mult_21_n364) );
  NOR2_X1 p6_mult_21_U520 ( .A1(p6_mult_21_n673), .A2(p6_mult_21_n708), .ZN(
        p6_mult_21_n365) );
  AOI21_X1 p6_mult_21_U519 ( .B1(p6_mult_21_n693), .B2(p6_mult_21_n691), .A(
        p6_mult_21_n707), .ZN(p6_mult_21_n706) );
  INV_X1 p6_mult_21_U518 ( .A(p6_mult_21_n706), .ZN(p6_mult_21_n366) );
  XNOR2_X1 p6_mult_21_U517 ( .A(B0[11]), .B(reg1_reg[7]), .ZN(p6_mult_21_n704)
         );
  OAI22_X1 p6_mult_21_U516 ( .A1(p6_mult_21_n704), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n705), .ZN(p6_mult_21_n367) );
  XNOR2_X1 p6_mult_21_U515 ( .A(B0[10]), .B(reg1_reg[7]), .ZN(p6_mult_21_n703)
         );
  OAI22_X1 p6_mult_21_U514 ( .A1(p6_mult_21_n703), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n704), .ZN(p6_mult_21_n368) );
  XNOR2_X1 p6_mult_21_U513 ( .A(B0[9]), .B(reg1_reg[7]), .ZN(p6_mult_21_n702)
         );
  OAI22_X1 p6_mult_21_U512 ( .A1(p6_mult_21_n702), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n703), .ZN(p6_mult_21_n369) );
  XNOR2_X1 p6_mult_21_U511 ( .A(B0[8]), .B(reg1_reg[7]), .ZN(p6_mult_21_n701)
         );
  OAI22_X1 p6_mult_21_U510 ( .A1(p6_mult_21_n701), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n702), .ZN(p6_mult_21_n370) );
  XNOR2_X1 p6_mult_21_U509 ( .A(B0[7]), .B(reg1_reg[7]), .ZN(p6_mult_21_n700)
         );
  OAI22_X1 p6_mult_21_U508 ( .A1(p6_mult_21_n700), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n701), .ZN(p6_mult_21_n371) );
  XNOR2_X1 p6_mult_21_U507 ( .A(B0[6]), .B(reg1_reg[7]), .ZN(p6_mult_21_n699)
         );
  OAI22_X1 p6_mult_21_U506 ( .A1(p6_mult_21_n699), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n700), .ZN(p6_mult_21_n372) );
  XNOR2_X1 p6_mult_21_U505 ( .A(B0[5]), .B(reg1_reg[7]), .ZN(p6_mult_21_n698)
         );
  OAI22_X1 p6_mult_21_U504 ( .A1(p6_mult_21_n698), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n699), .ZN(p6_mult_21_n373) );
  XNOR2_X1 p6_mult_21_U503 ( .A(B0[4]), .B(reg1_reg[7]), .ZN(p6_mult_21_n697)
         );
  OAI22_X1 p6_mult_21_U502 ( .A1(p6_mult_21_n697), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n698), .ZN(p6_mult_21_n374) );
  XNOR2_X1 p6_mult_21_U501 ( .A(B0[3]), .B(reg1_reg[7]), .ZN(p6_mult_21_n696)
         );
  OAI22_X1 p6_mult_21_U500 ( .A1(p6_mult_21_n696), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n697), .ZN(p6_mult_21_n375) );
  XNOR2_X1 p6_mult_21_U499 ( .A(B0[2]), .B(reg1_reg[7]), .ZN(p6_mult_21_n695)
         );
  OAI22_X1 p6_mult_21_U498 ( .A1(p6_mult_21_n695), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n696), .ZN(p6_mult_21_n376) );
  XNOR2_X1 p6_mult_21_U497 ( .A(B0[1]), .B(reg1_reg[7]), .ZN(p6_mult_21_n694)
         );
  OAI22_X1 p6_mult_21_U496 ( .A1(p6_mult_21_n694), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n695), .ZN(p6_mult_21_n377) );
  XNOR2_X1 p6_mult_21_U495 ( .A(reg1_reg[7]), .B(B0[0]), .ZN(p6_mult_21_n692)
         );
  OAI22_X1 p6_mult_21_U494 ( .A1(p6_mult_21_n692), .A2(p6_mult_21_n693), .B1(
        p6_mult_21_n691), .B2(p6_mult_21_n694), .ZN(p6_mult_21_n378) );
  NOR2_X1 p6_mult_21_U493 ( .A1(p6_mult_21_n673), .A2(p6_mult_21_n691), .ZN(
        p6_mult_21_n379) );
  AOI21_X1 p6_mult_21_U492 ( .B1(p6_mult_21_n676), .B2(p6_mult_21_n674), .A(
        p6_mult_21_n690), .ZN(p6_mult_21_n689) );
  INV_X1 p6_mult_21_U491 ( .A(p6_mult_21_n689), .ZN(p6_mult_21_n380) );
  XNOR2_X1 p6_mult_21_U490 ( .A(B0[11]), .B(reg1_reg[5]), .ZN(p6_mult_21_n687)
         );
  OAI22_X1 p6_mult_21_U489 ( .A1(p6_mult_21_n687), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n688), .ZN(p6_mult_21_n381) );
  OAI22_X1 p6_mult_21_U488 ( .A1(p6_mult_21_n686), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n687), .ZN(p6_mult_21_n382) );
  XNOR2_X1 p6_mult_21_U487 ( .A(B0[8]), .B(reg1_reg[5]), .ZN(p6_mult_21_n684)
         );
  OAI22_X1 p6_mult_21_U486 ( .A1(p6_mult_21_n684), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n685), .ZN(p6_mult_21_n384) );
  XNOR2_X1 p6_mult_21_U485 ( .A(B0[7]), .B(reg1_reg[5]), .ZN(p6_mult_21_n683)
         );
  OAI22_X1 p6_mult_21_U484 ( .A1(p6_mult_21_n683), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n684), .ZN(p6_mult_21_n385) );
  XNOR2_X1 p6_mult_21_U483 ( .A(B0[6]), .B(reg1_reg[5]), .ZN(p6_mult_21_n682)
         );
  OAI22_X1 p6_mult_21_U482 ( .A1(p6_mult_21_n682), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n683), .ZN(p6_mult_21_n386) );
  XNOR2_X1 p6_mult_21_U481 ( .A(B0[5]), .B(reg1_reg[5]), .ZN(p6_mult_21_n681)
         );
  OAI22_X1 p6_mult_21_U480 ( .A1(p6_mult_21_n681), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n682), .ZN(p6_mult_21_n387) );
  XNOR2_X1 p6_mult_21_U479 ( .A(B0[4]), .B(reg1_reg[5]), .ZN(p6_mult_21_n680)
         );
  OAI22_X1 p6_mult_21_U478 ( .A1(p6_mult_21_n680), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n681), .ZN(p6_mult_21_n388) );
  XNOR2_X1 p6_mult_21_U477 ( .A(B0[3]), .B(reg1_reg[5]), .ZN(p6_mult_21_n679)
         );
  OAI22_X1 p6_mult_21_U476 ( .A1(p6_mult_21_n679), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n680), .ZN(p6_mult_21_n389) );
  XNOR2_X1 p6_mult_21_U475 ( .A(B0[2]), .B(reg1_reg[5]), .ZN(p6_mult_21_n678)
         );
  OAI22_X1 p6_mult_21_U474 ( .A1(p6_mult_21_n678), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n679), .ZN(p6_mult_21_n390) );
  XNOR2_X1 p6_mult_21_U473 ( .A(B0[1]), .B(reg1_reg[5]), .ZN(p6_mult_21_n677)
         );
  OAI22_X1 p6_mult_21_U472 ( .A1(p6_mult_21_n677), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n678), .ZN(p6_mult_21_n391) );
  XNOR2_X1 p6_mult_21_U471 ( .A(reg1_reg[5]), .B(B0[0]), .ZN(p6_mult_21_n675)
         );
  OAI22_X1 p6_mult_21_U470 ( .A1(p6_mult_21_n675), .A2(p6_mult_21_n676), .B1(
        p6_mult_21_n674), .B2(p6_mult_21_n677), .ZN(p6_mult_21_n392) );
  NOR2_X1 p6_mult_21_U469 ( .A1(p6_mult_21_n673), .A2(p6_mult_21_n674), .ZN(
        p6_mult_21_n393) );
  AOI21_X1 p6_mult_21_U468 ( .B1(p6_mult_21_n657), .B2(p6_mult_21_n658), .A(
        p6_mult_21_n672), .ZN(p6_mult_21_n671) );
  INV_X1 p6_mult_21_U467 ( .A(p6_mult_21_n671), .ZN(p6_mult_21_n394) );
  XNOR2_X1 p6_mult_21_U466 ( .A(B0[11]), .B(reg1_reg[3]), .ZN(p6_mult_21_n669)
         );
  OAI22_X1 p6_mult_21_U465 ( .A1(p6_mult_21_n669), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n670), .ZN(p6_mult_21_n395) );
  XNOR2_X1 p6_mult_21_U464 ( .A(B0[10]), .B(reg1_reg[3]), .ZN(p6_mult_21_n668)
         );
  OAI22_X1 p6_mult_21_U463 ( .A1(p6_mult_21_n668), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n669), .ZN(p6_mult_21_n396) );
  XNOR2_X1 p6_mult_21_U462 ( .A(B0[9]), .B(reg1_reg[3]), .ZN(p6_mult_21_n667)
         );
  OAI22_X1 p6_mult_21_U461 ( .A1(p6_mult_21_n667), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n668), .ZN(p6_mult_21_n397) );
  XNOR2_X1 p6_mult_21_U460 ( .A(B0[8]), .B(reg1_reg[3]), .ZN(p6_mult_21_n666)
         );
  OAI22_X1 p6_mult_21_U459 ( .A1(p6_mult_21_n666), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n667), .ZN(p6_mult_21_n398) );
  XNOR2_X1 p6_mult_21_U458 ( .A(B0[7]), .B(reg1_reg[3]), .ZN(p6_mult_21_n665)
         );
  OAI22_X1 p6_mult_21_U457 ( .A1(p6_mult_21_n665), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n666), .ZN(p6_mult_21_n399) );
  XNOR2_X1 p6_mult_21_U456 ( .A(B0[6]), .B(reg1_reg[3]), .ZN(p6_mult_21_n664)
         );
  OAI22_X1 p6_mult_21_U455 ( .A1(p6_mult_21_n664), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n665), .ZN(p6_mult_21_n400) );
  XNOR2_X1 p6_mult_21_U454 ( .A(B0[5]), .B(reg1_reg[3]), .ZN(p6_mult_21_n663)
         );
  OAI22_X1 p6_mult_21_U453 ( .A1(p6_mult_21_n663), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n664), .ZN(p6_mult_21_n401) );
  XNOR2_X1 p6_mult_21_U452 ( .A(B0[4]), .B(reg1_reg[3]), .ZN(p6_mult_21_n662)
         );
  OAI22_X1 p6_mult_21_U451 ( .A1(p6_mult_21_n662), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n663), .ZN(p6_mult_21_n402) );
  XNOR2_X1 p6_mult_21_U450 ( .A(B0[3]), .B(reg1_reg[3]), .ZN(p6_mult_21_n661)
         );
  OAI22_X1 p6_mult_21_U449 ( .A1(p6_mult_21_n661), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n662), .ZN(p6_mult_21_n403) );
  XNOR2_X1 p6_mult_21_U448 ( .A(B0[2]), .B(reg1_reg[3]), .ZN(p6_mult_21_n660)
         );
  OAI22_X1 p6_mult_21_U447 ( .A1(p6_mult_21_n660), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n661), .ZN(p6_mult_21_n404) );
  XNOR2_X1 p6_mult_21_U446 ( .A(B0[1]), .B(reg1_reg[3]), .ZN(p6_mult_21_n659)
         );
  OAI22_X1 p6_mult_21_U445 ( .A1(p6_mult_21_n659), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n660), .ZN(p6_mult_21_n405) );
  XNOR2_X1 p6_mult_21_U444 ( .A(reg1_reg[3]), .B(B0[0]), .ZN(p6_mult_21_n656)
         );
  OAI22_X1 p6_mult_21_U443 ( .A1(p6_mult_21_n656), .A2(p6_mult_21_n657), .B1(
        p6_mult_21_n658), .B2(p6_mult_21_n659), .ZN(p6_mult_21_n406) );
  XOR2_X1 p6_mult_21_U442 ( .A(B0[13]), .B(p6_mult_21_n655), .Z(
        p6_mult_21_n653) );
  AOI21_X1 p6_mult_21_U441 ( .B1(p6_mult_21_n641), .B2(p6_mult_21_n643), .A(
        p6_mult_21_n653), .ZN(p6_mult_21_n654) );
  INV_X1 p6_mult_21_U440 ( .A(p6_mult_21_n654), .ZN(p6_mult_21_n408) );
  XNOR2_X1 p6_mult_21_U439 ( .A(B0[12]), .B(reg1_reg[1]), .ZN(p6_mult_21_n652)
         );
  OAI22_X1 p6_mult_21_U438 ( .A1(p6_mult_21_n652), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n653), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n409) );
  XNOR2_X1 p6_mult_21_U437 ( .A(B0[11]), .B(reg1_reg[1]), .ZN(p6_mult_21_n651)
         );
  OAI22_X1 p6_mult_21_U436 ( .A1(p6_mult_21_n651), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n652), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n410) );
  XNOR2_X1 p6_mult_21_U435 ( .A(B0[10]), .B(reg1_reg[1]), .ZN(p6_mult_21_n650)
         );
  OAI22_X1 p6_mult_21_U434 ( .A1(p6_mult_21_n650), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n651), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n411) );
  XNOR2_X1 p6_mult_21_U433 ( .A(B0[9]), .B(reg1_reg[1]), .ZN(p6_mult_21_n649)
         );
  OAI22_X1 p6_mult_21_U432 ( .A1(p6_mult_21_n649), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n650), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n412) );
  XNOR2_X1 p6_mult_21_U431 ( .A(B0[8]), .B(reg1_reg[1]), .ZN(p6_mult_21_n648)
         );
  OAI22_X1 p6_mult_21_U430 ( .A1(p6_mult_21_n648), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n649), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n413) );
  XNOR2_X1 p6_mult_21_U429 ( .A(B0[7]), .B(reg1_reg[1]), .ZN(p6_mult_21_n647)
         );
  OAI22_X1 p6_mult_21_U428 ( .A1(p6_mult_21_n647), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n648), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n414) );
  XNOR2_X1 p6_mult_21_U427 ( .A(B0[6]), .B(reg1_reg[1]), .ZN(p6_mult_21_n646)
         );
  OAI22_X1 p6_mult_21_U426 ( .A1(p6_mult_21_n646), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n647), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n415) );
  XNOR2_X1 p6_mult_21_U425 ( .A(B0[5]), .B(reg1_reg[1]), .ZN(p6_mult_21_n645)
         );
  OAI22_X1 p6_mult_21_U424 ( .A1(p6_mult_21_n645), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n646), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n416) );
  XNOR2_X1 p6_mult_21_U423 ( .A(B0[4]), .B(reg1_reg[1]), .ZN(p6_mult_21_n644)
         );
  OAI22_X1 p6_mult_21_U422 ( .A1(p6_mult_21_n644), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n645), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n417) );
  XNOR2_X1 p6_mult_21_U421 ( .A(B0[3]), .B(reg1_reg[1]), .ZN(p6_mult_21_n642)
         );
  OAI22_X1 p6_mult_21_U420 ( .A1(p6_mult_21_n642), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n644), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n418) );
  OAI22_X1 p6_mult_21_U419 ( .A1(p6_mult_21_n640), .A2(p6_mult_21_n641), .B1(
        p6_mult_21_n642), .B2(p6_mult_21_n643), .ZN(p6_mult_21_n419) );
  OAI21_X1 p6_mult_21_U418 ( .B1(p6_mult_21_n637), .B2(p6_mult_21_n638), .A(
        p6_mult_21_n639), .ZN(p6_mult_21_n636) );
  XOR2_X1 p6_mult_21_U417 ( .A(p6_mult_21_n636), .B(p6_mult_21_n136), .Z(
        p6_mult_21_n635) );
  XNOR2_X1 p6_mult_21_U416 ( .A(p6_mult_21_n162), .B(p6_mult_21_n635), .ZN(
        temp1[13]) );
  XOR2_X2 p6_mult_21_U415 ( .A(reg1_reg[12]), .B(p6_mult_21_n764), .Z(
        p6_mult_21_n742) );
  XOR2_X2 p6_mult_21_U414 ( .A(reg1_reg[10]), .B(p6_mult_21_n762), .Z(
        p6_mult_21_n725) );
  XOR2_X2 p6_mult_21_U413 ( .A(reg1_reg[8]), .B(p6_mult_21_n760), .Z(
        p6_mult_21_n708) );
  XOR2_X2 p6_mult_21_U412 ( .A(reg1_reg[6]), .B(p6_mult_21_n758), .Z(
        p6_mult_21_n691) );
  XOR2_X2 p6_mult_21_U411 ( .A(reg1_reg[4]), .B(p6_mult_21_n771), .Z(
        p6_mult_21_n674) );
  INV_X1 p6_mult_21_U410 ( .A(reg1_reg[0]), .ZN(p6_mult_21_n643) );
  INV_X1 p6_mult_21_U409 ( .A(p6_mult_21_n798), .ZN(p6_mult_21_n658) );
  HA_X1 p6_mult_21_U145 ( .A(p6_mult_21_n406), .B(p6_mult_21_n419), .CO(
        p6_mult_21_n315), .S(p6_mult_21_n316) );
  FA_X1 p6_mult_21_U144 ( .A(p6_mult_21_n418), .B(p6_mult_21_n393), .CI(
        p6_mult_21_n405), .CO(p6_mult_21_n313), .S(p6_mult_21_n314) );
  HA_X1 p6_mult_21_U143 ( .A(p6_mult_21_n321), .B(p6_mult_21_n392), .CO(
        p6_mult_21_n311), .S(p6_mult_21_n312) );
  FA_X1 p6_mult_21_U142 ( .A(p6_mult_21_n404), .B(p6_mult_21_n417), .CI(
        p6_mult_21_n312), .CO(p6_mult_21_n309), .S(p6_mult_21_n310) );
  FA_X1 p6_mult_21_U141 ( .A(p6_mult_21_n416), .B(p6_mult_21_n379), .CI(
        p6_mult_21_n403), .CO(p6_mult_21_n307), .S(p6_mult_21_n308) );
  FA_X1 p6_mult_21_U140 ( .A(p6_mult_21_n311), .B(p6_mult_21_n391), .CI(
        p6_mult_21_n308), .CO(p6_mult_21_n305), .S(p6_mult_21_n306) );
  HA_X1 p6_mult_21_U139 ( .A(p6_mult_21_n320), .B(p6_mult_21_n378), .CO(
        p6_mult_21_n303), .S(p6_mult_21_n304) );
  FA_X1 p6_mult_21_U138 ( .A(p6_mult_21_n390), .B(p6_mult_21_n415), .CI(
        p6_mult_21_n402), .CO(p6_mult_21_n301), .S(p6_mult_21_n302) );
  FA_X1 p6_mult_21_U137 ( .A(p6_mult_21_n307), .B(p6_mult_21_n304), .CI(
        p6_mult_21_n302), .CO(p6_mult_21_n299), .S(p6_mult_21_n300) );
  FA_X1 p6_mult_21_U136 ( .A(p6_mult_21_n389), .B(p6_mult_21_n365), .CI(
        p6_mult_21_n414), .CO(p6_mult_21_n297), .S(p6_mult_21_n298) );
  FA_X1 p6_mult_21_U135 ( .A(p6_mult_21_n377), .B(p6_mult_21_n401), .CI(
        p6_mult_21_n303), .CO(p6_mult_21_n295), .S(p6_mult_21_n296) );
  FA_X1 p6_mult_21_U134 ( .A(p6_mult_21_n298), .B(p6_mult_21_n301), .CI(
        p6_mult_21_n296), .CO(p6_mult_21_n293), .S(p6_mult_21_n294) );
  HA_X1 p6_mult_21_U133 ( .A(p6_mult_21_n319), .B(p6_mult_21_n364), .CO(
        p6_mult_21_n291), .S(p6_mult_21_n292) );
  FA_X1 p6_mult_21_U132 ( .A(p6_mult_21_n376), .B(p6_mult_21_n388), .CI(
        p6_mult_21_n400), .CO(p6_mult_21_n289), .S(p6_mult_21_n290) );
  FA_X1 p6_mult_21_U131 ( .A(p6_mult_21_n292), .B(p6_mult_21_n413), .CI(
        p6_mult_21_n297), .CO(p6_mult_21_n287), .S(p6_mult_21_n288) );
  FA_X1 p6_mult_21_U130 ( .A(p6_mult_21_n290), .B(p6_mult_21_n295), .CI(
        p6_mult_21_n288), .CO(p6_mult_21_n285), .S(p6_mult_21_n286) );
  FA_X1 p6_mult_21_U129 ( .A(p6_mult_21_n375), .B(p6_mult_21_n351), .CI(
        p6_mult_21_n412), .CO(p6_mult_21_n283), .S(p6_mult_21_n284) );
  FA_X1 p6_mult_21_U128 ( .A(p6_mult_21_n363), .B(p6_mult_21_n399), .CI(
        p6_mult_21_n387), .CO(p6_mult_21_n281), .S(p6_mult_21_n282) );
  FA_X1 p6_mult_21_U127 ( .A(p6_mult_21_n289), .B(p6_mult_21_n291), .CI(
        p6_mult_21_n284), .CO(p6_mult_21_n279), .S(p6_mult_21_n280) );
  FA_X1 p6_mult_21_U126 ( .A(p6_mult_21_n287), .B(p6_mult_21_n282), .CI(
        p6_mult_21_n280), .CO(p6_mult_21_n277), .S(p6_mult_21_n278) );
  HA_X1 p6_mult_21_U125 ( .A(p6_mult_21_n318), .B(p6_mult_21_n350), .CO(
        p6_mult_21_n275), .S(p6_mult_21_n276) );
  FA_X1 p6_mult_21_U124 ( .A(p6_mult_21_n362), .B(p6_mult_21_n386), .CI(
        p6_mult_21_n411), .CO(p6_mult_21_n273), .S(p6_mult_21_n274) );
  FA_X1 p6_mult_21_U123 ( .A(p6_mult_21_n374), .B(p6_mult_21_n398), .CI(
        p6_mult_21_n276), .CO(p6_mult_21_n271), .S(p6_mult_21_n272) );
  FA_X1 p6_mult_21_U122 ( .A(p6_mult_21_n281), .B(p6_mult_21_n283), .CI(
        p6_mult_21_n274), .CO(p6_mult_21_n269), .S(p6_mult_21_n270) );
  FA_X1 p6_mult_21_U121 ( .A(p6_mult_21_n279), .B(p6_mult_21_n272), .CI(
        p6_mult_21_n270), .CO(p6_mult_21_n267), .S(p6_mult_21_n268) );
  FA_X1 p6_mult_21_U120 ( .A(p6_mult_21_n361), .B(p6_mult_21_n337), .CI(
        p6_mult_21_n410), .CO(p6_mult_21_n265), .S(p6_mult_21_n266) );
  FA_X1 p6_mult_21_U109 ( .A(p6_mult_21_n349), .B(p6_mult_21_n397), .CI(
        p6_mult_21_n373), .CO(p6_mult_21_n263), .S(p6_mult_21_n264) );
  FA_X1 p6_mult_21_U108 ( .A(p6_mult_21_n275), .B(p6_mult_21_n385), .CI(
        p6_mult_21_n273), .CO(p6_mult_21_n261), .S(p6_mult_21_n262) );
  FA_X1 p6_mult_21_U107 ( .A(p6_mult_21_n264), .B(p6_mult_21_n266), .CI(
        p6_mult_21_n271), .CO(p6_mult_21_n259), .S(p6_mult_21_n260) );
  FA_X1 p6_mult_21_U106 ( .A(p6_mult_21_n262), .B(p6_mult_21_n269), .CI(
        p6_mult_21_n260), .CO(p6_mult_21_n257), .S(p6_mult_21_n258) );
  HA_X1 p6_mult_21_U105 ( .A(p6_mult_21_n317), .B(p6_mult_21_n336), .CO(
        p6_mult_21_n255), .S(p6_mult_21_n256) );
  FA_X1 p6_mult_21_U104 ( .A(p6_mult_21_n409), .B(p6_mult_21_n372), .CI(
        p6_mult_21_n396), .CO(p6_mult_21_n253), .S(p6_mult_21_n254) );
  FA_X1 p6_mult_21_U103 ( .A(p6_mult_21_n348), .B(p6_mult_21_n384), .CI(
        p6_mult_21_n360), .CO(p6_mult_21_n251), .S(p6_mult_21_n252) );
  FA_X1 p6_mult_21_U102 ( .A(p6_mult_21_n265), .B(p6_mult_21_n256), .CI(
        p6_mult_21_n263), .CO(p6_mult_21_n249), .S(p6_mult_21_n250) );
  FA_X1 p6_mult_21_U101 ( .A(p6_mult_21_n254), .B(p6_mult_21_n252), .CI(
        p6_mult_21_n261), .CO(p6_mult_21_n247), .S(p6_mult_21_n248) );
  FA_X1 p6_mult_21_U100 ( .A(p6_mult_21_n259), .B(p6_mult_21_n250), .CI(
        p6_mult_21_n248), .CO(p6_mult_21_n245), .S(p6_mult_21_n246) );
  FA_X1 p6_mult_21_U97 ( .A(p6_mult_21_n395), .B(p6_mult_21_n359), .CI(
        p6_mult_21_n408), .CO(p6_mult_21_n241), .S(p6_mult_21_n242) );
  FA_X1 p6_mult_21_U96 ( .A(p6_mult_21_n335), .B(p6_mult_21_n371), .CI(
        p6_mult_21_n255), .CO(p6_mult_21_n239), .S(p6_mult_21_n240) );
  FA_X1 p6_mult_21_U95 ( .A(p6_mult_21_n253), .B(p6_mult_21_n244), .CI(
        p6_mult_21_n251), .CO(p6_mult_21_n237), .S(p6_mult_21_n238) );
  FA_X1 p6_mult_21_U94 ( .A(p6_mult_21_n240), .B(p6_mult_21_n242), .CI(
        p6_mult_21_n249), .CO(p6_mult_21_n235), .S(p6_mult_21_n236) );
  FA_X1 p6_mult_21_U93 ( .A(p6_mult_21_n247), .B(p6_mult_21_n238), .CI(
        p6_mult_21_n236), .CO(p6_mult_21_n233), .S(p6_mult_21_n234) );
  FA_X1 p6_mult_21_U91 ( .A(p6_mult_21_n382), .B(p6_mult_21_n346), .CI(
        p6_mult_21_n232), .CO(p6_mult_21_n229), .S(p6_mult_21_n230) );
  FA_X1 p6_mult_21_U90 ( .A(p6_mult_21_n334), .B(p6_mult_21_n370), .CI(
        p6_mult_21_n358), .CO(p6_mult_21_n227), .S(p6_mult_21_n228) );
  FA_X1 p6_mult_21_U89 ( .A(p6_mult_21_n241), .B(p6_mult_21_n243), .CI(
        p6_mult_21_n239), .CO(p6_mult_21_n225), .S(p6_mult_21_n226) );
  FA_X1 p6_mult_21_U88 ( .A(p6_mult_21_n230), .B(p6_mult_21_n228), .CI(
        p6_mult_21_n237), .CO(p6_mult_21_n223), .S(p6_mult_21_n224) );
  FA_X1 p6_mult_21_U87 ( .A(p6_mult_21_n235), .B(p6_mult_21_n226), .CI(
        p6_mult_21_n224), .CO(p6_mult_21_n221), .S(p6_mult_21_n222) );
  FA_X1 p6_mult_21_U86 ( .A(p6_mult_21_n231), .B(p6_mult_21_n333), .CI(
        p6_mult_21_n394), .CO(p6_mult_21_n219), .S(p6_mult_21_n220) );
  FA_X1 p6_mult_21_U85 ( .A(p6_mult_21_n345), .B(p6_mult_21_n381), .CI(
        p6_mult_21_n357), .CO(p6_mult_21_n217), .S(p6_mult_21_n218) );
  FA_X1 p6_mult_21_U84 ( .A(p6_mult_21_n229), .B(p6_mult_21_n369), .CI(
        p6_mult_21_n227), .CO(p6_mult_21_n215), .S(p6_mult_21_n216) );
  FA_X1 p6_mult_21_U83 ( .A(p6_mult_21_n220), .B(p6_mult_21_n218), .CI(
        p6_mult_21_n225), .CO(p6_mult_21_n213), .S(p6_mult_21_n214) );
  FA_X1 p6_mult_21_U82 ( .A(p6_mult_21_n223), .B(p6_mult_21_n216), .CI(
        p6_mult_21_n214), .CO(p6_mult_21_n211), .S(p6_mult_21_n212) );
  FA_X1 p6_mult_21_U80 ( .A(p6_mult_21_n368), .B(p6_mult_21_n344), .CI(
        p6_mult_21_n210), .CO(p6_mult_21_n207), .S(p6_mult_21_n208) );
  FA_X1 p6_mult_21_U79 ( .A(p6_mult_21_n332), .B(p6_mult_21_n356), .CI(
        p6_mult_21_n219), .CO(p6_mult_21_n205), .S(p6_mult_21_n206) );
  FA_X1 p6_mult_21_U78 ( .A(p6_mult_21_n208), .B(p6_mult_21_n217), .CI(
        p6_mult_21_n215), .CO(p6_mult_21_n203), .S(p6_mult_21_n204) );
  FA_X1 p6_mult_21_U77 ( .A(p6_mult_21_n213), .B(p6_mult_21_n206), .CI(
        p6_mult_21_n204), .CO(p6_mult_21_n201), .S(p6_mult_21_n202) );
  FA_X1 p6_mult_21_U76 ( .A(p6_mult_21_n209), .B(p6_mult_21_n331), .CI(
        p6_mult_21_n380), .CO(p6_mult_21_n199), .S(p6_mult_21_n200) );
  FA_X1 p6_mult_21_U75 ( .A(p6_mult_21_n355), .B(p6_mult_21_n343), .CI(
        p6_mult_21_n367), .CO(p6_mult_21_n197), .S(p6_mult_21_n198) );
  FA_X1 p6_mult_21_U74 ( .A(p6_mult_21_n198), .B(p6_mult_21_n207), .CI(
        p6_mult_21_n200), .CO(p6_mult_21_n195), .S(p6_mult_21_n196) );
  FA_X1 p6_mult_21_U73 ( .A(p6_mult_21_n203), .B(p6_mult_21_n205), .CI(
        p6_mult_21_n196), .CO(p6_mult_21_n193), .S(p6_mult_21_n194) );
  FA_X1 p6_mult_21_U71 ( .A(p6_mult_21_n330), .B(p6_mult_21_n342), .CI(
        p6_mult_21_n192), .CO(p6_mult_21_n189), .S(p6_mult_21_n190) );
  FA_X1 p6_mult_21_U70 ( .A(p6_mult_21_n199), .B(p6_mult_21_n354), .CI(
        p6_mult_21_n197), .CO(p6_mult_21_n187), .S(p6_mult_21_n188) );
  FA_X1 p6_mult_21_U69 ( .A(p6_mult_21_n188), .B(p6_mult_21_n190), .CI(
        p6_mult_21_n195), .CO(p6_mult_21_n185), .S(p6_mult_21_n186) );
  FA_X1 p6_mult_21_U68 ( .A(p6_mult_21_n191), .B(p6_mult_21_n329), .CI(
        p6_mult_21_n366), .CO(p6_mult_21_n183), .S(p6_mult_21_n184) );
  FA_X1 p6_mult_21_U67 ( .A(p6_mult_21_n341), .B(p6_mult_21_n353), .CI(
        p6_mult_21_n189), .CO(p6_mult_21_n181), .S(p6_mult_21_n182) );
  FA_X1 p6_mult_21_U66 ( .A(p6_mult_21_n187), .B(p6_mult_21_n184), .CI(
        p6_mult_21_n182), .CO(p6_mult_21_n179), .S(p6_mult_21_n180) );
  FA_X1 p6_mult_21_U64 ( .A(p6_mult_21_n328), .B(p6_mult_21_n340), .CI(
        p6_mult_21_n178), .CO(p6_mult_21_n175), .S(p6_mult_21_n176) );
  FA_X1 p6_mult_21_U63 ( .A(p6_mult_21_n176), .B(p6_mult_21_n183), .CI(
        p6_mult_21_n181), .CO(p6_mult_21_n173), .S(p6_mult_21_n174) );
  FA_X1 p6_mult_21_U62 ( .A(p6_mult_21_n327), .B(p6_mult_21_n177), .CI(
        p6_mult_21_n352), .CO(p6_mult_21_n171), .S(p6_mult_21_n172) );
  FA_X1 p6_mult_21_U61 ( .A(p6_mult_21_n175), .B(p6_mult_21_n339), .CI(
        p6_mult_21_n172), .CO(p6_mult_21_n169), .S(p6_mult_21_n170) );
  FA_X1 p6_mult_21_U59 ( .A(p6_mult_21_n168), .B(p6_mult_21_n326), .CI(
        p6_mult_21_n171), .CO(p6_mult_21_n165), .S(p6_mult_21_n166) );
  FA_X1 p6_mult_21_U58 ( .A(p6_mult_21_n325), .B(p6_mult_21_n167), .CI(
        p6_mult_21_n338), .CO(p6_mult_21_n163), .S(p6_mult_21_n164) );
  FA_X1 p6_mult_21_U44 ( .A(p6_mult_21_n246), .B(p6_mult_21_n257), .CI(
        p6_mult_21_n149), .CO(p6_mult_21_n148), .S(temp1[0]) );
  FA_X1 p6_mult_21_U43 ( .A(p6_mult_21_n234), .B(p6_mult_21_n245), .CI(
        p6_mult_21_n148), .CO(p6_mult_21_n147), .S(temp1[1]) );
  FA_X1 p6_mult_21_U42 ( .A(p6_mult_21_n222), .B(p6_mult_21_n233), .CI(
        p6_mult_21_n147), .CO(p6_mult_21_n146), .S(temp1[2]) );
  FA_X1 p6_mult_21_U41 ( .A(p6_mult_21_n212), .B(p6_mult_21_n221), .CI(
        p6_mult_21_n146), .CO(p6_mult_21_n145), .S(temp1[3]) );
  FA_X1 p6_mult_21_U40 ( .A(p6_mult_21_n202), .B(p6_mult_21_n211), .CI(
        p6_mult_21_n145), .CO(p6_mult_21_n144), .S(temp1[4]) );
  FA_X1 p6_mult_21_U39 ( .A(p6_mult_21_n194), .B(p6_mult_21_n201), .CI(
        p6_mult_21_n144), .CO(p6_mult_21_n143), .S(temp1[5]) );
  FA_X1 p6_mult_21_U38 ( .A(p6_mult_21_n186), .B(p6_mult_21_n193), .CI(
        p6_mult_21_n143), .CO(p6_mult_21_n142), .S(temp1[6]) );
  FA_X1 p6_mult_21_U37 ( .A(p6_mult_21_n180), .B(p6_mult_21_n185), .CI(
        p6_mult_21_n142), .CO(p6_mult_21_n141), .S(temp1[7]) );
  FA_X1 p6_mult_21_U30 ( .A(p6_mult_21_n174), .B(p6_mult_21_n179), .CI(
        p6_mult_21_n141), .CO(p6_mult_21_n140), .S(temp1[8]) );
  FA_X1 p6_mult_21_U20 ( .A(p6_mult_21_n170), .B(p6_mult_21_n173), .CI(
        p6_mult_21_n140), .CO(p6_mult_21_n139), .S(temp1[9]) );
  FA_X1 p6_mult_21_U10 ( .A(p6_mult_21_n166), .B(p6_mult_21_n169), .CI(
        p6_mult_21_n139), .CO(p6_mult_21_n138), .S(temp1[10]) );
  FA_X1 p6_mult_21_U9 ( .A(p6_mult_21_n165), .B(p6_mult_21_n164), .CI(
        p6_mult_21_n138), .CO(p6_mult_21_n137), .S(temp1[11]) );
  FA_X1 p6_mult_21_U8 ( .A(p6_mult_21_n163), .B(p6_mult_21_n162), .CI(
        p6_mult_21_n137), .CO(p6_mult_21_n136), .S(temp1[12]) );
  NAND2_X1 REG1_1_U34 ( .A1(temp1[4]), .A2(REG1_1_n43), .ZN(REG1_1_n85) );
  OAI21_X1 REG1_1_U33 ( .B1(REG1_1_n45), .B2(REG1_1_n66), .A(REG1_1_n85), .ZN(
        REG1_1_n57) );
  NAND2_X1 REG1_1_U32 ( .A1(temp1[3]), .A2(REG1_1_n43), .ZN(REG1_1_n86) );
  OAI21_X1 REG1_1_U31 ( .B1(REG1_1_n45), .B2(REG1_1_n65), .A(REG1_1_n86), .ZN(
        REG1_1_n58) );
  NAND2_X1 REG1_1_U30 ( .A1(temp1[2]), .A2(REG1_1_n43), .ZN(REG1_1_n87) );
  OAI21_X1 REG1_1_U29 ( .B1(REG1_1_n45), .B2(REG1_1_n64), .A(REG1_1_n87), .ZN(
        REG1_1_n59) );
  NAND2_X1 REG1_1_U28 ( .A1(temp1[5]), .A2(REG1_1_n43), .ZN(REG1_1_n84) );
  OAI21_X1 REG1_1_U27 ( .B1(REG1_1_n44), .B2(REG1_1_n67), .A(REG1_1_n84), .ZN(
        REG1_1_n56) );
  NAND2_X1 REG1_1_U26 ( .A1(temp1[9]), .A2(REG1_1_n43), .ZN(REG1_1_n80) );
  OAI21_X1 REG1_1_U25 ( .B1(REG1_1_n44), .B2(REG1_1_n71), .A(REG1_1_n80), .ZN(
        REG1_1_n52) );
  NAND2_X1 REG1_1_U24 ( .A1(temp1[8]), .A2(REG1_1_n44), .ZN(REG1_1_n81) );
  OAI21_X1 REG1_1_U23 ( .B1(REG1_1_n44), .B2(REG1_1_n70), .A(REG1_1_n81), .ZN(
        REG1_1_n53) );
  NAND2_X1 REG1_1_U22 ( .A1(temp1[7]), .A2(REG1_1_n43), .ZN(REG1_1_n82) );
  OAI21_X1 REG1_1_U21 ( .B1(REG1_1_n44), .B2(REG1_1_n69), .A(REG1_1_n82), .ZN(
        REG1_1_n54) );
  NAND2_X1 REG1_1_U20 ( .A1(temp1[6]), .A2(REG1_1_n43), .ZN(REG1_1_n83) );
  OAI21_X1 REG1_1_U19 ( .B1(REG1_1_n44), .B2(REG1_1_n68), .A(REG1_1_n83), .ZN(
        REG1_1_n55) );
  NAND2_X1 REG1_1_U18 ( .A1(temp1[1]), .A2(REG1_1_n43), .ZN(REG1_1_n88) );
  OAI21_X1 REG1_1_U17 ( .B1(REG1_1_n44), .B2(REG1_1_n63), .A(REG1_1_n88), .ZN(
        REG1_1_n60) );
  NAND2_X1 REG1_1_U16 ( .A1(temp1[0]), .A2(REG1_1_n43), .ZN(REG1_1_n89) );
  OAI21_X1 REG1_1_U15 ( .B1(REG1_1_n44), .B2(REG1_1_n62), .A(REG1_1_n89), .ZN(
        REG1_1_n61) );
  NAND2_X1 REG1_1_U14 ( .A1(temp1[10]), .A2(REG1_1_n44), .ZN(REG1_1_n79) );
  OAI21_X1 REG1_1_U13 ( .B1(REG1_1_n44), .B2(REG1_1_n72), .A(REG1_1_n79), .ZN(
        REG1_1_n51) );
  NAND2_X1 REG1_1_U12 ( .A1(temp1[12]), .A2(REG1_1_n43), .ZN(REG1_1_n77) );
  OAI21_X1 REG1_1_U11 ( .B1(REG1_1_n44), .B2(REG1_1_n74), .A(REG1_1_n77), .ZN(
        REG1_1_n49) );
  NAND2_X1 REG1_1_U10 ( .A1(temp1[11]), .A2(REG1_1_n43), .ZN(REG1_1_n78) );
  OAI21_X1 REG1_1_U9 ( .B1(REG1_1_n44), .B2(REG1_1_n73), .A(REG1_1_n78), .ZN(
        REG1_1_n50) );
  NAND2_X1 REG1_1_U8 ( .A1(temp1[13]), .A2(REG1_1_n43), .ZN(REG1_1_n76) );
  OAI21_X1 REG1_1_U7 ( .B1(REG1_1_n44), .B2(REG1_1_n75), .A(REG1_1_n76), .ZN(
        REG1_1_n48) );
  BUF_X1 REG1_1_U6 ( .A(n47), .Z(REG1_1_n47) );
  BUF_X1 REG1_1_U5 ( .A(n47), .Z(REG1_1_n46) );
  BUF_X1 REG1_1_U4 ( .A(VIN), .Z(REG1_1_n45) );
  BUF_X1 REG1_1_U3 ( .A(VIN), .Z(REG1_1_n43) );
  BUF_X1 REG1_1_U2 ( .A(VIN), .Z(REG1_1_n44) );
  DFFR_X1 REG1_1_q_reg_0_ ( .D(REG1_1_n61), .CK(CLK), .RN(REG1_1_n47), .Q(
        mul1_reg[0]), .QN(REG1_1_n62) );
  DFFR_X1 REG1_1_q_reg_1_ ( .D(REG1_1_n60), .CK(CLK), .RN(REG1_1_n47), .Q(
        mul1_reg[1]), .QN(REG1_1_n63) );
  DFFR_X1 REG1_1_q_reg_2_ ( .D(REG1_1_n59), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[2]), .QN(REG1_1_n64) );
  DFFR_X1 REG1_1_q_reg_3_ ( .D(REG1_1_n58), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[3]), .QN(REG1_1_n65) );
  DFFR_X1 REG1_1_q_reg_4_ ( .D(REG1_1_n57), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[4]), .QN(REG1_1_n66) );
  DFFR_X1 REG1_1_q_reg_5_ ( .D(REG1_1_n56), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[5]), .QN(REG1_1_n67) );
  DFFR_X1 REG1_1_q_reg_6_ ( .D(REG1_1_n55), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[6]), .QN(REG1_1_n68) );
  DFFR_X1 REG1_1_q_reg_7_ ( .D(REG1_1_n54), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[7]), .QN(REG1_1_n69) );
  DFFR_X1 REG1_1_q_reg_8_ ( .D(REG1_1_n53), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[8]), .QN(REG1_1_n70) );
  DFFR_X1 REG1_1_q_reg_9_ ( .D(REG1_1_n52), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[9]), .QN(REG1_1_n71) );
  DFFR_X1 REG1_1_q_reg_10_ ( .D(REG1_1_n51), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[10]), .QN(REG1_1_n72) );
  DFFR_X1 REG1_1_q_reg_11_ ( .D(REG1_1_n50), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[11]), .QN(REG1_1_n73) );
  DFFR_X1 REG1_1_q_reg_12_ ( .D(REG1_1_n49), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[12]), .QN(REG1_1_n74) );
  DFFR_X1 REG1_1_q_reg_13_ ( .D(REG1_1_n48), .CK(CLK), .RN(REG1_1_n46), .Q(
        mul1_reg[13]), .QN(REG1_1_n75) );
  NAND2_X1 REGISTER2_U34 ( .A1(reg2[3]), .A2(REGISTER2_n43), .ZN(REGISTER2_n86) );
  OAI21_X1 REGISTER2_U33 ( .B1(REGISTER2_n45), .B2(REGISTER2_n65), .A(
        REGISTER2_n86), .ZN(REGISTER2_n58) );
  NAND2_X1 REGISTER2_U32 ( .A1(reg2[12]), .A2(REGISTER2_n43), .ZN(
        REGISTER2_n77) );
  OAI21_X1 REGISTER2_U31 ( .B1(REGISTER2_n44), .B2(REGISTER2_n74), .A(
        REGISTER2_n77), .ZN(REGISTER2_n49) );
  NAND2_X1 REGISTER2_U30 ( .A1(reg2[6]), .A2(REGISTER2_n43), .ZN(REGISTER2_n83) );
  OAI21_X1 REGISTER2_U29 ( .B1(REGISTER2_n44), .B2(REGISTER2_n68), .A(
        REGISTER2_n83), .ZN(REGISTER2_n55) );
  NAND2_X1 REGISTER2_U28 ( .A1(reg2[4]), .A2(REGISTER2_n43), .ZN(REGISTER2_n85) );
  OAI21_X1 REGISTER2_U27 ( .B1(REGISTER2_n45), .B2(REGISTER2_n66), .A(
        REGISTER2_n85), .ZN(REGISTER2_n57) );
  NAND2_X1 REGISTER2_U26 ( .A1(reg2[2]), .A2(REGISTER2_n43), .ZN(REGISTER2_n87) );
  OAI21_X1 REGISTER2_U25 ( .B1(REGISTER2_n45), .B2(REGISTER2_n64), .A(
        REGISTER2_n87), .ZN(REGISTER2_n59) );
  NAND2_X1 REGISTER2_U24 ( .A1(reg2[0]), .A2(REGISTER2_n43), .ZN(REGISTER2_n89) );
  OAI21_X1 REGISTER2_U23 ( .B1(REGISTER2_n44), .B2(REGISTER2_n62), .A(
        REGISTER2_n89), .ZN(REGISTER2_n61) );
  NAND2_X1 REGISTER2_U22 ( .A1(reg2[13]), .A2(REGISTER2_n43), .ZN(
        REGISTER2_n76) );
  OAI21_X1 REGISTER2_U21 ( .B1(REGISTER2_n44), .B2(REGISTER2_n75), .A(
        REGISTER2_n76), .ZN(REGISTER2_n48) );
  NAND2_X1 REGISTER2_U20 ( .A1(reg2[10]), .A2(REGISTER2_n44), .ZN(
        REGISTER2_n79) );
  OAI21_X1 REGISTER2_U19 ( .B1(REGISTER2_n44), .B2(REGISTER2_n72), .A(
        REGISTER2_n79), .ZN(REGISTER2_n51) );
  NAND2_X1 REGISTER2_U18 ( .A1(reg2[8]), .A2(REGISTER2_n44), .ZN(REGISTER2_n81) );
  OAI21_X1 REGISTER2_U17 ( .B1(REGISTER2_n44), .B2(REGISTER2_n70), .A(
        REGISTER2_n81), .ZN(REGISTER2_n53) );
  NAND2_X1 REGISTER2_U16 ( .A1(reg2[1]), .A2(REGISTER2_n43), .ZN(REGISTER2_n88) );
  OAI21_X1 REGISTER2_U15 ( .B1(REGISTER2_n44), .B2(REGISTER2_n63), .A(
        REGISTER2_n88), .ZN(REGISTER2_n60) );
  NAND2_X1 REGISTER2_U14 ( .A1(reg2[11]), .A2(REGISTER2_n43), .ZN(
        REGISTER2_n78) );
  OAI21_X1 REGISTER2_U13 ( .B1(REGISTER2_n44), .B2(REGISTER2_n73), .A(
        REGISTER2_n78), .ZN(REGISTER2_n50) );
  NAND2_X1 REGISTER2_U12 ( .A1(reg2[9]), .A2(REGISTER2_n43), .ZN(REGISTER2_n80) );
  OAI21_X1 REGISTER2_U11 ( .B1(REGISTER2_n44), .B2(REGISTER2_n71), .A(
        REGISTER2_n80), .ZN(REGISTER2_n52) );
  NAND2_X1 REGISTER2_U10 ( .A1(reg2[7]), .A2(REGISTER2_n43), .ZN(REGISTER2_n82) );
  OAI21_X1 REGISTER2_U9 ( .B1(REGISTER2_n44), .B2(REGISTER2_n69), .A(
        REGISTER2_n82), .ZN(REGISTER2_n54) );
  NAND2_X1 REGISTER2_U8 ( .A1(reg2[5]), .A2(REGISTER2_n43), .ZN(REGISTER2_n84)
         );
  OAI21_X1 REGISTER2_U7 ( .B1(REGISTER2_n44), .B2(REGISTER2_n67), .A(
        REGISTER2_n84), .ZN(REGISTER2_n56) );
  BUF_X1 REGISTER2_U6 ( .A(n47), .Z(REGISTER2_n47) );
  BUF_X1 REGISTER2_U5 ( .A(n47), .Z(REGISTER2_n46) );
  BUF_X1 REGISTER2_U4 ( .A(VIN), .Z(REGISTER2_n45) );
  BUF_X1 REGISTER2_U3 ( .A(VIN), .Z(REGISTER2_n43) );
  BUF_X1 REGISTER2_U2 ( .A(VIN), .Z(REGISTER2_n44) );
  DFFR_X1 REGISTER2_q_reg_0_ ( .D(REGISTER2_n61), .CK(CLK), .RN(REGISTER2_n47), 
        .Q(reg2_reg[0]), .QN(REGISTER2_n62) );
  DFFR_X1 REGISTER2_q_reg_1_ ( .D(REGISTER2_n60), .CK(CLK), .RN(REGISTER2_n47), 
        .Q(reg2_reg[1]), .QN(REGISTER2_n63) );
  DFFR_X1 REGISTER2_q_reg_2_ ( .D(REGISTER2_n59), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[2]), .QN(REGISTER2_n64) );
  DFFR_X1 REGISTER2_q_reg_3_ ( .D(REGISTER2_n58), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[3]), .QN(REGISTER2_n65) );
  DFFR_X1 REGISTER2_q_reg_4_ ( .D(REGISTER2_n57), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[4]), .QN(REGISTER2_n66) );
  DFFR_X1 REGISTER2_q_reg_5_ ( .D(REGISTER2_n56), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[5]), .QN(REGISTER2_n67) );
  DFFR_X1 REGISTER2_q_reg_6_ ( .D(REGISTER2_n55), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[6]), .QN(REGISTER2_n68) );
  DFFR_X1 REGISTER2_q_reg_7_ ( .D(REGISTER2_n54), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[7]), .QN(REGISTER2_n69) );
  DFFR_X1 REGISTER2_q_reg_8_ ( .D(REGISTER2_n53), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[8]), .QN(REGISTER2_n70) );
  DFFR_X1 REGISTER2_q_reg_9_ ( .D(REGISTER2_n52), .CK(CLK), .RN(REGISTER2_n46), 
        .Q(reg2_reg[9]), .QN(REGISTER2_n71) );
  DFFR_X1 REGISTER2_q_reg_10_ ( .D(REGISTER2_n51), .CK(CLK), .RN(REGISTER2_n46), .Q(reg2_reg[10]), .QN(REGISTER2_n72) );
  DFFR_X1 REGISTER2_q_reg_11_ ( .D(REGISTER2_n50), .CK(CLK), .RN(REGISTER2_n46), .Q(reg2_reg[11]), .QN(REGISTER2_n73) );
  DFFR_X1 REGISTER2_q_reg_12_ ( .D(REGISTER2_n49), .CK(CLK), .RN(REGISTER2_n46), .Q(reg2_reg[12]), .QN(REGISTER2_n74) );
  DFFR_X1 REGISTER2_q_reg_13_ ( .D(REGISTER2_n48), .CK(CLK), .RN(REGISTER2_n46), .Q(reg2_reg[13]), .QN(REGISTER2_n75) );
  XOR2_X1 p7_mult_21_U691 ( .A(reg2_reg[2]), .B(reg2_reg[1]), .Z(
        p7_mult_21_n798) );
  INV_X1 p7_mult_21_U690 ( .A(reg2_reg[1]), .ZN(p7_mult_21_n655) );
  NOR2_X1 p7_mult_21_U689 ( .A1(p7_mult_21_n655), .A2(B1[1]), .ZN(
        p7_mult_21_n803) );
  INV_X1 p7_mult_21_U688 ( .A(p7_mult_21_n803), .ZN(p7_mult_21_n805) );
  NAND2_X1 p7_mult_21_U687 ( .A1(reg2_reg[1]), .A2(p7_mult_21_n643), .ZN(
        p7_mult_21_n641) );
  XNOR2_X1 p7_mult_21_U686 ( .A(B1[2]), .B(reg2_reg[1]), .ZN(p7_mult_21_n640)
         );
  OAI22_X1 p7_mult_21_U685 ( .A1(p7_mult_21_n805), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n640), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n804) );
  NAND2_X1 p7_mult_21_U684 ( .A1(p7_mult_21_n798), .A2(p7_mult_21_n804), .ZN(
        p7_mult_21_n801) );
  NAND2_X1 p7_mult_21_U683 ( .A1(p7_mult_21_n803), .A2(p7_mult_21_n804), .ZN(
        p7_mult_21_n802) );
  INV_X1 p7_mult_21_U682 ( .A(B1[0]), .ZN(p7_mult_21_n673) );
  MUX2_X1 p7_mult_21_U681 ( .A(p7_mult_21_n801), .B(p7_mult_21_n802), .S(
        p7_mult_21_n673), .Z(p7_mult_21_n800) );
  INV_X1 p7_mult_21_U680 ( .A(p7_mult_21_n800), .ZN(p7_mult_21_n795) );
  INV_X1 p7_mult_21_U679 ( .A(reg2_reg[3]), .ZN(p7_mult_21_n771) );
  XNOR2_X1 p7_mult_21_U678 ( .A(p7_mult_21_n771), .B(reg2_reg[2]), .ZN(
        p7_mult_21_n799) );
  NAND2_X1 p7_mult_21_U677 ( .A1(p7_mult_21_n658), .A2(p7_mult_21_n799), .ZN(
        p7_mult_21_n657) );
  NAND3_X1 p7_mult_21_U676 ( .A1(p7_mult_21_n798), .A2(p7_mult_21_n673), .A3(
        reg2_reg[3]), .ZN(p7_mult_21_n797) );
  OAI21_X1 p7_mult_21_U675 ( .B1(p7_mult_21_n771), .B2(p7_mult_21_n657), .A(
        p7_mult_21_n797), .ZN(p7_mult_21_n796) );
  AOI222_X1 p7_mult_21_U674 ( .A1(p7_mult_21_n795), .A2(p7_mult_21_n316), .B1(
        p7_mult_21_n796), .B2(p7_mult_21_n795), .C1(p7_mult_21_n796), .C2(
        p7_mult_21_n316), .ZN(p7_mult_21_n794) );
  INV_X1 p7_mult_21_U673 ( .A(p7_mult_21_n794), .ZN(p7_mult_21_n793) );
  AOI222_X1 p7_mult_21_U672 ( .A1(p7_mult_21_n793), .A2(p7_mult_21_n314), .B1(
        p7_mult_21_n793), .B2(p7_mult_21_n315), .C1(p7_mult_21_n315), .C2(
        p7_mult_21_n314), .ZN(p7_mult_21_n792) );
  INV_X1 p7_mult_21_U671 ( .A(p7_mult_21_n792), .ZN(p7_mult_21_n791) );
  AOI222_X1 p7_mult_21_U670 ( .A1(p7_mult_21_n791), .A2(p7_mult_21_n310), .B1(
        p7_mult_21_n791), .B2(p7_mult_21_n313), .C1(p7_mult_21_n313), .C2(
        p7_mult_21_n310), .ZN(p7_mult_21_n790) );
  INV_X1 p7_mult_21_U669 ( .A(p7_mult_21_n790), .ZN(p7_mult_21_n789) );
  AOI222_X1 p7_mult_21_U668 ( .A1(p7_mult_21_n789), .A2(p7_mult_21_n306), .B1(
        p7_mult_21_n789), .B2(p7_mult_21_n309), .C1(p7_mult_21_n309), .C2(
        p7_mult_21_n306), .ZN(p7_mult_21_n788) );
  INV_X1 p7_mult_21_U667 ( .A(p7_mult_21_n788), .ZN(p7_mult_21_n787) );
  AOI222_X1 p7_mult_21_U666 ( .A1(p7_mult_21_n787), .A2(p7_mult_21_n300), .B1(
        p7_mult_21_n787), .B2(p7_mult_21_n305), .C1(p7_mult_21_n305), .C2(
        p7_mult_21_n300), .ZN(p7_mult_21_n786) );
  INV_X1 p7_mult_21_U665 ( .A(p7_mult_21_n786), .ZN(p7_mult_21_n785) );
  AOI222_X1 p7_mult_21_U664 ( .A1(p7_mult_21_n785), .A2(p7_mult_21_n294), .B1(
        p7_mult_21_n785), .B2(p7_mult_21_n299), .C1(p7_mult_21_n299), .C2(
        p7_mult_21_n294), .ZN(p7_mult_21_n784) );
  INV_X1 p7_mult_21_U663 ( .A(p7_mult_21_n784), .ZN(p7_mult_21_n783) );
  AOI222_X1 p7_mult_21_U662 ( .A1(p7_mult_21_n783), .A2(p7_mult_21_n286), .B1(
        p7_mult_21_n783), .B2(p7_mult_21_n293), .C1(p7_mult_21_n293), .C2(
        p7_mult_21_n286), .ZN(p7_mult_21_n780) );
  INV_X1 p7_mult_21_U661 ( .A(p7_mult_21_n278), .ZN(p7_mult_21_n781) );
  INV_X1 p7_mult_21_U660 ( .A(p7_mult_21_n285), .ZN(p7_mult_21_n782) );
  OAI222_X1 p7_mult_21_U659 ( .A1(p7_mult_21_n780), .A2(p7_mult_21_n781), .B1(
        p7_mult_21_n780), .B2(p7_mult_21_n782), .C1(p7_mult_21_n782), .C2(
        p7_mult_21_n781), .ZN(p7_mult_21_n779) );
  AOI222_X1 p7_mult_21_U658 ( .A1(p7_mult_21_n779), .A2(p7_mult_21_n268), .B1(
        p7_mult_21_n779), .B2(p7_mult_21_n277), .C1(p7_mult_21_n277), .C2(
        p7_mult_21_n268), .ZN(p7_mult_21_n776) );
  INV_X1 p7_mult_21_U657 ( .A(p7_mult_21_n258), .ZN(p7_mult_21_n777) );
  INV_X1 p7_mult_21_U656 ( .A(p7_mult_21_n267), .ZN(p7_mult_21_n778) );
  OAI222_X1 p7_mult_21_U655 ( .A1(p7_mult_21_n776), .A2(p7_mult_21_n777), .B1(
        p7_mult_21_n776), .B2(p7_mult_21_n778), .C1(p7_mult_21_n778), .C2(
        p7_mult_21_n777), .ZN(p7_mult_21_n149) );
  XOR2_X1 p7_mult_21_U654 ( .A(B1[12]), .B(reg2_reg[13]), .Z(p7_mult_21_n757)
         );
  INV_X1 p7_mult_21_U653 ( .A(reg2_reg[11]), .ZN(p7_mult_21_n764) );
  INV_X1 p7_mult_21_U652 ( .A(reg2_reg[13]), .ZN(p7_mult_21_n766) );
  XNOR2_X1 p7_mult_21_U651 ( .A(p7_mult_21_n766), .B(reg2_reg[12]), .ZN(
        p7_mult_21_n775) );
  NAND2_X1 p7_mult_21_U650 ( .A1(p7_mult_21_n742), .A2(p7_mult_21_n775), .ZN(
        p7_mult_21_n744) );
  INV_X1 p7_mult_21_U649 ( .A(p7_mult_21_n744), .ZN(p7_mult_21_n637) );
  INV_X1 p7_mult_21_U648 ( .A(p7_mult_21_n742), .ZN(p7_mult_21_n638) );
  XNOR2_X1 p7_mult_21_U647 ( .A(B1[13]), .B(p7_mult_21_n766), .ZN(
        p7_mult_21_n639) );
  AOI22_X1 p7_mult_21_U646 ( .A1(p7_mult_21_n757), .A2(p7_mult_21_n637), .B1(
        p7_mult_21_n638), .B2(p7_mult_21_n639), .ZN(p7_mult_21_n162) );
  XNOR2_X1 p7_mult_21_U645 ( .A(B1[12]), .B(reg2_reg[11]), .ZN(p7_mult_21_n739) );
  INV_X1 p7_mult_21_U644 ( .A(reg2_reg[9]), .ZN(p7_mult_21_n762) );
  XNOR2_X1 p7_mult_21_U643 ( .A(p7_mult_21_n764), .B(reg2_reg[10]), .ZN(
        p7_mult_21_n774) );
  NAND2_X1 p7_mult_21_U642 ( .A1(p7_mult_21_n725), .A2(p7_mult_21_n774), .ZN(
        p7_mult_21_n727) );
  XNOR2_X1 p7_mult_21_U641 ( .A(B1[13]), .B(reg2_reg[11]), .ZN(p7_mult_21_n741) );
  OAI22_X1 p7_mult_21_U640 ( .A1(p7_mult_21_n739), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n741), .ZN(p7_mult_21_n167) );
  INV_X1 p7_mult_21_U639 ( .A(p7_mult_21_n167), .ZN(p7_mult_21_n168) );
  XNOR2_X1 p7_mult_21_U638 ( .A(B1[12]), .B(reg2_reg[9]), .ZN(p7_mult_21_n722)
         );
  INV_X1 p7_mult_21_U637 ( .A(reg2_reg[7]), .ZN(p7_mult_21_n760) );
  XNOR2_X1 p7_mult_21_U636 ( .A(p7_mult_21_n762), .B(reg2_reg[8]), .ZN(
        p7_mult_21_n773) );
  NAND2_X1 p7_mult_21_U635 ( .A1(p7_mult_21_n708), .A2(p7_mult_21_n773), .ZN(
        p7_mult_21_n710) );
  XNOR2_X1 p7_mult_21_U634 ( .A(B1[13]), .B(reg2_reg[9]), .ZN(p7_mult_21_n724)
         );
  OAI22_X1 p7_mult_21_U633 ( .A1(p7_mult_21_n722), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n724), .ZN(p7_mult_21_n177) );
  INV_X1 p7_mult_21_U632 ( .A(p7_mult_21_n177), .ZN(p7_mult_21_n178) );
  XNOR2_X1 p7_mult_21_U631 ( .A(B1[12]), .B(reg2_reg[7]), .ZN(p7_mult_21_n705)
         );
  INV_X1 p7_mult_21_U630 ( .A(reg2_reg[5]), .ZN(p7_mult_21_n758) );
  XNOR2_X1 p7_mult_21_U629 ( .A(p7_mult_21_n760), .B(reg2_reg[6]), .ZN(
        p7_mult_21_n772) );
  NAND2_X1 p7_mult_21_U628 ( .A1(p7_mult_21_n691), .A2(p7_mult_21_n772), .ZN(
        p7_mult_21_n693) );
  XNOR2_X1 p7_mult_21_U627 ( .A(B1[13]), .B(reg2_reg[7]), .ZN(p7_mult_21_n707)
         );
  OAI22_X1 p7_mult_21_U626 ( .A1(p7_mult_21_n705), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n707), .ZN(p7_mult_21_n191) );
  INV_X1 p7_mult_21_U625 ( .A(p7_mult_21_n191), .ZN(p7_mult_21_n192) );
  XNOR2_X1 p7_mult_21_U624 ( .A(B1[12]), .B(reg2_reg[5]), .ZN(p7_mult_21_n688)
         );
  XNOR2_X1 p7_mult_21_U623 ( .A(p7_mult_21_n758), .B(reg2_reg[4]), .ZN(
        p7_mult_21_n770) );
  NAND2_X1 p7_mult_21_U622 ( .A1(p7_mult_21_n674), .A2(p7_mult_21_n770), .ZN(
        p7_mult_21_n676) );
  XNOR2_X1 p7_mult_21_U621 ( .A(B1[13]), .B(reg2_reg[5]), .ZN(p7_mult_21_n690)
         );
  OAI22_X1 p7_mult_21_U620 ( .A1(p7_mult_21_n688), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n690), .ZN(p7_mult_21_n209) );
  INV_X1 p7_mult_21_U619 ( .A(p7_mult_21_n209), .ZN(p7_mult_21_n210) );
  XNOR2_X1 p7_mult_21_U618 ( .A(B1[12]), .B(reg2_reg[3]), .ZN(p7_mult_21_n670)
         );
  XNOR2_X1 p7_mult_21_U617 ( .A(B1[13]), .B(reg2_reg[3]), .ZN(p7_mult_21_n672)
         );
  OAI22_X1 p7_mult_21_U616 ( .A1(p7_mult_21_n670), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n672), .ZN(p7_mult_21_n231) );
  INV_X1 p7_mult_21_U615 ( .A(p7_mult_21_n231), .ZN(p7_mult_21_n232) );
  XNOR2_X1 p7_mult_21_U614 ( .A(B1[3]), .B(reg2_reg[11]), .ZN(p7_mult_21_n730)
         );
  XNOR2_X1 p7_mult_21_U613 ( .A(B1[4]), .B(reg2_reg[11]), .ZN(p7_mult_21_n731)
         );
  OAI22_X1 p7_mult_21_U612 ( .A1(p7_mult_21_n730), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n731), .ZN(p7_mult_21_n768) );
  XNOR2_X1 p7_mult_21_U611 ( .A(B1[9]), .B(reg2_reg[5]), .ZN(p7_mult_21_n685)
         );
  XNOR2_X1 p7_mult_21_U610 ( .A(B1[10]), .B(reg2_reg[5]), .ZN(p7_mult_21_n686)
         );
  OAI22_X1 p7_mult_21_U609 ( .A1(p7_mult_21_n685), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n686), .ZN(p7_mult_21_n769) );
  OR2_X1 p7_mult_21_U608 ( .A1(p7_mult_21_n768), .A2(p7_mult_21_n769), .ZN(
        p7_mult_21_n243) );
  XNOR2_X1 p7_mult_21_U607 ( .A(p7_mult_21_n768), .B(p7_mult_21_n769), .ZN(
        p7_mult_21_n244) );
  NAND3_X1 p7_mult_21_U606 ( .A1(p7_mult_21_n638), .A2(p7_mult_21_n673), .A3(
        reg2_reg[13]), .ZN(p7_mult_21_n767) );
  OAI21_X1 p7_mult_21_U605 ( .B1(p7_mult_21_n766), .B2(p7_mult_21_n744), .A(
        p7_mult_21_n767), .ZN(p7_mult_21_n317) );
  OR3_X1 p7_mult_21_U604 ( .A1(p7_mult_21_n725), .A2(B1[0]), .A3(
        p7_mult_21_n764), .ZN(p7_mult_21_n765) );
  OAI21_X1 p7_mult_21_U603 ( .B1(p7_mult_21_n764), .B2(p7_mult_21_n727), .A(
        p7_mult_21_n765), .ZN(p7_mult_21_n318) );
  OR3_X1 p7_mult_21_U602 ( .A1(p7_mult_21_n708), .A2(B1[0]), .A3(
        p7_mult_21_n762), .ZN(p7_mult_21_n763) );
  OAI21_X1 p7_mult_21_U601 ( .B1(p7_mult_21_n762), .B2(p7_mult_21_n710), .A(
        p7_mult_21_n763), .ZN(p7_mult_21_n319) );
  OR3_X1 p7_mult_21_U600 ( .A1(p7_mult_21_n691), .A2(B1[0]), .A3(
        p7_mult_21_n760), .ZN(p7_mult_21_n761) );
  OAI21_X1 p7_mult_21_U599 ( .B1(p7_mult_21_n760), .B2(p7_mult_21_n693), .A(
        p7_mult_21_n761), .ZN(p7_mult_21_n320) );
  OR3_X1 p7_mult_21_U598 ( .A1(p7_mult_21_n674), .A2(B1[0]), .A3(
        p7_mult_21_n758), .ZN(p7_mult_21_n759) );
  OAI21_X1 p7_mult_21_U597 ( .B1(p7_mult_21_n758), .B2(p7_mult_21_n676), .A(
        p7_mult_21_n759), .ZN(p7_mult_21_n321) );
  XNOR2_X1 p7_mult_21_U596 ( .A(B1[11]), .B(reg2_reg[13]), .ZN(p7_mult_21_n755) );
  INV_X1 p7_mult_21_U595 ( .A(p7_mult_21_n757), .ZN(p7_mult_21_n756) );
  OAI22_X1 p7_mult_21_U594 ( .A1(p7_mult_21_n755), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n756), .ZN(p7_mult_21_n325) );
  XNOR2_X1 p7_mult_21_U593 ( .A(B1[10]), .B(reg2_reg[13]), .ZN(p7_mult_21_n754) );
  OAI22_X1 p7_mult_21_U592 ( .A1(p7_mult_21_n754), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n755), .ZN(p7_mult_21_n326) );
  XNOR2_X1 p7_mult_21_U591 ( .A(B1[9]), .B(reg2_reg[13]), .ZN(p7_mult_21_n753)
         );
  OAI22_X1 p7_mult_21_U590 ( .A1(p7_mult_21_n753), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n754), .ZN(p7_mult_21_n327) );
  XNOR2_X1 p7_mult_21_U589 ( .A(B1[8]), .B(reg2_reg[13]), .ZN(p7_mult_21_n752)
         );
  OAI22_X1 p7_mult_21_U588 ( .A1(p7_mult_21_n752), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n753), .ZN(p7_mult_21_n328) );
  XNOR2_X1 p7_mult_21_U587 ( .A(B1[7]), .B(reg2_reg[13]), .ZN(p7_mult_21_n751)
         );
  OAI22_X1 p7_mult_21_U586 ( .A1(p7_mult_21_n751), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n752), .ZN(p7_mult_21_n329) );
  XNOR2_X1 p7_mult_21_U585 ( .A(B1[6]), .B(reg2_reg[13]), .ZN(p7_mult_21_n750)
         );
  OAI22_X1 p7_mult_21_U584 ( .A1(p7_mult_21_n750), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n751), .ZN(p7_mult_21_n330) );
  XNOR2_X1 p7_mult_21_U583 ( .A(B1[5]), .B(reg2_reg[13]), .ZN(p7_mult_21_n749)
         );
  OAI22_X1 p7_mult_21_U582 ( .A1(p7_mult_21_n749), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n750), .ZN(p7_mult_21_n331) );
  XNOR2_X1 p7_mult_21_U581 ( .A(B1[4]), .B(reg2_reg[13]), .ZN(p7_mult_21_n748)
         );
  OAI22_X1 p7_mult_21_U580 ( .A1(p7_mult_21_n748), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n749), .ZN(p7_mult_21_n332) );
  XNOR2_X1 p7_mult_21_U579 ( .A(B1[3]), .B(reg2_reg[13]), .ZN(p7_mult_21_n747)
         );
  OAI22_X1 p7_mult_21_U578 ( .A1(p7_mult_21_n747), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n748), .ZN(p7_mult_21_n333) );
  XNOR2_X1 p7_mult_21_U577 ( .A(B1[2]), .B(reg2_reg[13]), .ZN(p7_mult_21_n746)
         );
  OAI22_X1 p7_mult_21_U576 ( .A1(p7_mult_21_n746), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n747), .ZN(p7_mult_21_n334) );
  XNOR2_X1 p7_mult_21_U575 ( .A(B1[1]), .B(reg2_reg[13]), .ZN(p7_mult_21_n745)
         );
  OAI22_X1 p7_mult_21_U574 ( .A1(p7_mult_21_n745), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n746), .ZN(p7_mult_21_n335) );
  XNOR2_X1 p7_mult_21_U573 ( .A(reg2_reg[13]), .B(B1[0]), .ZN(p7_mult_21_n743)
         );
  OAI22_X1 p7_mult_21_U572 ( .A1(p7_mult_21_n743), .A2(p7_mult_21_n744), .B1(
        p7_mult_21_n742), .B2(p7_mult_21_n745), .ZN(p7_mult_21_n336) );
  NOR2_X1 p7_mult_21_U571 ( .A1(p7_mult_21_n673), .A2(p7_mult_21_n742), .ZN(
        p7_mult_21_n337) );
  AOI21_X1 p7_mult_21_U570 ( .B1(p7_mult_21_n727), .B2(p7_mult_21_n725), .A(
        p7_mult_21_n741), .ZN(p7_mult_21_n740) );
  INV_X1 p7_mult_21_U569 ( .A(p7_mult_21_n740), .ZN(p7_mult_21_n338) );
  XNOR2_X1 p7_mult_21_U568 ( .A(B1[11]), .B(reg2_reg[11]), .ZN(p7_mult_21_n738) );
  OAI22_X1 p7_mult_21_U567 ( .A1(p7_mult_21_n738), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n739), .ZN(p7_mult_21_n339) );
  XNOR2_X1 p7_mult_21_U566 ( .A(B1[10]), .B(reg2_reg[11]), .ZN(p7_mult_21_n737) );
  OAI22_X1 p7_mult_21_U565 ( .A1(p7_mult_21_n737), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n738), .ZN(p7_mult_21_n340) );
  XNOR2_X1 p7_mult_21_U564 ( .A(B1[9]), .B(reg2_reg[11]), .ZN(p7_mult_21_n736)
         );
  OAI22_X1 p7_mult_21_U563 ( .A1(p7_mult_21_n736), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n737), .ZN(p7_mult_21_n341) );
  XNOR2_X1 p7_mult_21_U562 ( .A(B1[8]), .B(reg2_reg[11]), .ZN(p7_mult_21_n735)
         );
  OAI22_X1 p7_mult_21_U561 ( .A1(p7_mult_21_n735), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n736), .ZN(p7_mult_21_n342) );
  XNOR2_X1 p7_mult_21_U560 ( .A(B1[7]), .B(reg2_reg[11]), .ZN(p7_mult_21_n734)
         );
  OAI22_X1 p7_mult_21_U559 ( .A1(p7_mult_21_n734), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n735), .ZN(p7_mult_21_n343) );
  XNOR2_X1 p7_mult_21_U558 ( .A(B1[6]), .B(reg2_reg[11]), .ZN(p7_mult_21_n733)
         );
  OAI22_X1 p7_mult_21_U557 ( .A1(p7_mult_21_n733), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n734), .ZN(p7_mult_21_n344) );
  XNOR2_X1 p7_mult_21_U556 ( .A(B1[5]), .B(reg2_reg[11]), .ZN(p7_mult_21_n732)
         );
  OAI22_X1 p7_mult_21_U555 ( .A1(p7_mult_21_n732), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n733), .ZN(p7_mult_21_n345) );
  OAI22_X1 p7_mult_21_U554 ( .A1(p7_mult_21_n731), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n732), .ZN(p7_mult_21_n346) );
  XNOR2_X1 p7_mult_21_U553 ( .A(B1[2]), .B(reg2_reg[11]), .ZN(p7_mult_21_n729)
         );
  OAI22_X1 p7_mult_21_U552 ( .A1(p7_mult_21_n729), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n730), .ZN(p7_mult_21_n348) );
  XNOR2_X1 p7_mult_21_U551 ( .A(B1[1]), .B(reg2_reg[11]), .ZN(p7_mult_21_n728)
         );
  OAI22_X1 p7_mult_21_U550 ( .A1(p7_mult_21_n728), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n729), .ZN(p7_mult_21_n349) );
  XNOR2_X1 p7_mult_21_U549 ( .A(reg2_reg[11]), .B(B1[0]), .ZN(p7_mult_21_n726)
         );
  OAI22_X1 p7_mult_21_U548 ( .A1(p7_mult_21_n726), .A2(p7_mult_21_n727), .B1(
        p7_mult_21_n725), .B2(p7_mult_21_n728), .ZN(p7_mult_21_n350) );
  NOR2_X1 p7_mult_21_U547 ( .A1(p7_mult_21_n673), .A2(p7_mult_21_n725), .ZN(
        p7_mult_21_n351) );
  AOI21_X1 p7_mult_21_U546 ( .B1(p7_mult_21_n710), .B2(p7_mult_21_n708), .A(
        p7_mult_21_n724), .ZN(p7_mult_21_n723) );
  INV_X1 p7_mult_21_U545 ( .A(p7_mult_21_n723), .ZN(p7_mult_21_n352) );
  XNOR2_X1 p7_mult_21_U544 ( .A(B1[11]), .B(reg2_reg[9]), .ZN(p7_mult_21_n721)
         );
  OAI22_X1 p7_mult_21_U543 ( .A1(p7_mult_21_n721), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n722), .ZN(p7_mult_21_n353) );
  XNOR2_X1 p7_mult_21_U542 ( .A(B1[10]), .B(reg2_reg[9]), .ZN(p7_mult_21_n720)
         );
  OAI22_X1 p7_mult_21_U541 ( .A1(p7_mult_21_n720), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n721), .ZN(p7_mult_21_n354) );
  XNOR2_X1 p7_mult_21_U540 ( .A(B1[9]), .B(reg2_reg[9]), .ZN(p7_mult_21_n719)
         );
  OAI22_X1 p7_mult_21_U539 ( .A1(p7_mult_21_n719), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n720), .ZN(p7_mult_21_n355) );
  XNOR2_X1 p7_mult_21_U538 ( .A(B1[8]), .B(reg2_reg[9]), .ZN(p7_mult_21_n718)
         );
  OAI22_X1 p7_mult_21_U537 ( .A1(p7_mult_21_n718), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n719), .ZN(p7_mult_21_n356) );
  XNOR2_X1 p7_mult_21_U536 ( .A(B1[7]), .B(reg2_reg[9]), .ZN(p7_mult_21_n717)
         );
  OAI22_X1 p7_mult_21_U535 ( .A1(p7_mult_21_n717), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n718), .ZN(p7_mult_21_n357) );
  XNOR2_X1 p7_mult_21_U534 ( .A(B1[6]), .B(reg2_reg[9]), .ZN(p7_mult_21_n716)
         );
  OAI22_X1 p7_mult_21_U533 ( .A1(p7_mult_21_n716), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n717), .ZN(p7_mult_21_n358) );
  XNOR2_X1 p7_mult_21_U532 ( .A(B1[5]), .B(reg2_reg[9]), .ZN(p7_mult_21_n715)
         );
  OAI22_X1 p7_mult_21_U531 ( .A1(p7_mult_21_n715), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n716), .ZN(p7_mult_21_n359) );
  XNOR2_X1 p7_mult_21_U530 ( .A(B1[4]), .B(reg2_reg[9]), .ZN(p7_mult_21_n714)
         );
  OAI22_X1 p7_mult_21_U529 ( .A1(p7_mult_21_n714), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n715), .ZN(p7_mult_21_n360) );
  XNOR2_X1 p7_mult_21_U528 ( .A(B1[3]), .B(reg2_reg[9]), .ZN(p7_mult_21_n713)
         );
  OAI22_X1 p7_mult_21_U527 ( .A1(p7_mult_21_n713), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n714), .ZN(p7_mult_21_n361) );
  XNOR2_X1 p7_mult_21_U526 ( .A(B1[2]), .B(reg2_reg[9]), .ZN(p7_mult_21_n712)
         );
  OAI22_X1 p7_mult_21_U525 ( .A1(p7_mult_21_n712), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n713), .ZN(p7_mult_21_n362) );
  XNOR2_X1 p7_mult_21_U524 ( .A(B1[1]), .B(reg2_reg[9]), .ZN(p7_mult_21_n711)
         );
  OAI22_X1 p7_mult_21_U523 ( .A1(p7_mult_21_n711), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n712), .ZN(p7_mult_21_n363) );
  XNOR2_X1 p7_mult_21_U522 ( .A(reg2_reg[9]), .B(B1[0]), .ZN(p7_mult_21_n709)
         );
  OAI22_X1 p7_mult_21_U521 ( .A1(p7_mult_21_n709), .A2(p7_mult_21_n710), .B1(
        p7_mult_21_n708), .B2(p7_mult_21_n711), .ZN(p7_mult_21_n364) );
  NOR2_X1 p7_mult_21_U520 ( .A1(p7_mult_21_n673), .A2(p7_mult_21_n708), .ZN(
        p7_mult_21_n365) );
  AOI21_X1 p7_mult_21_U519 ( .B1(p7_mult_21_n693), .B2(p7_mult_21_n691), .A(
        p7_mult_21_n707), .ZN(p7_mult_21_n706) );
  INV_X1 p7_mult_21_U518 ( .A(p7_mult_21_n706), .ZN(p7_mult_21_n366) );
  XNOR2_X1 p7_mult_21_U517 ( .A(B1[11]), .B(reg2_reg[7]), .ZN(p7_mult_21_n704)
         );
  OAI22_X1 p7_mult_21_U516 ( .A1(p7_mult_21_n704), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n705), .ZN(p7_mult_21_n367) );
  XNOR2_X1 p7_mult_21_U515 ( .A(B1[10]), .B(reg2_reg[7]), .ZN(p7_mult_21_n703)
         );
  OAI22_X1 p7_mult_21_U514 ( .A1(p7_mult_21_n703), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n704), .ZN(p7_mult_21_n368) );
  XNOR2_X1 p7_mult_21_U513 ( .A(B1[9]), .B(reg2_reg[7]), .ZN(p7_mult_21_n702)
         );
  OAI22_X1 p7_mult_21_U512 ( .A1(p7_mult_21_n702), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n703), .ZN(p7_mult_21_n369) );
  XNOR2_X1 p7_mult_21_U511 ( .A(B1[8]), .B(reg2_reg[7]), .ZN(p7_mult_21_n701)
         );
  OAI22_X1 p7_mult_21_U510 ( .A1(p7_mult_21_n701), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n702), .ZN(p7_mult_21_n370) );
  XNOR2_X1 p7_mult_21_U509 ( .A(B1[7]), .B(reg2_reg[7]), .ZN(p7_mult_21_n700)
         );
  OAI22_X1 p7_mult_21_U508 ( .A1(p7_mult_21_n700), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n701), .ZN(p7_mult_21_n371) );
  XNOR2_X1 p7_mult_21_U507 ( .A(B1[6]), .B(reg2_reg[7]), .ZN(p7_mult_21_n699)
         );
  OAI22_X1 p7_mult_21_U506 ( .A1(p7_mult_21_n699), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n700), .ZN(p7_mult_21_n372) );
  XNOR2_X1 p7_mult_21_U505 ( .A(B1[5]), .B(reg2_reg[7]), .ZN(p7_mult_21_n698)
         );
  OAI22_X1 p7_mult_21_U504 ( .A1(p7_mult_21_n698), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n699), .ZN(p7_mult_21_n373) );
  XNOR2_X1 p7_mult_21_U503 ( .A(B1[4]), .B(reg2_reg[7]), .ZN(p7_mult_21_n697)
         );
  OAI22_X1 p7_mult_21_U502 ( .A1(p7_mult_21_n697), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n698), .ZN(p7_mult_21_n374) );
  XNOR2_X1 p7_mult_21_U501 ( .A(B1[3]), .B(reg2_reg[7]), .ZN(p7_mult_21_n696)
         );
  OAI22_X1 p7_mult_21_U500 ( .A1(p7_mult_21_n696), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n697), .ZN(p7_mult_21_n375) );
  XNOR2_X1 p7_mult_21_U499 ( .A(B1[2]), .B(reg2_reg[7]), .ZN(p7_mult_21_n695)
         );
  OAI22_X1 p7_mult_21_U498 ( .A1(p7_mult_21_n695), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n696), .ZN(p7_mult_21_n376) );
  XNOR2_X1 p7_mult_21_U497 ( .A(B1[1]), .B(reg2_reg[7]), .ZN(p7_mult_21_n694)
         );
  OAI22_X1 p7_mult_21_U496 ( .A1(p7_mult_21_n694), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n695), .ZN(p7_mult_21_n377) );
  XNOR2_X1 p7_mult_21_U495 ( .A(reg2_reg[7]), .B(B1[0]), .ZN(p7_mult_21_n692)
         );
  OAI22_X1 p7_mult_21_U494 ( .A1(p7_mult_21_n692), .A2(p7_mult_21_n693), .B1(
        p7_mult_21_n691), .B2(p7_mult_21_n694), .ZN(p7_mult_21_n378) );
  NOR2_X1 p7_mult_21_U493 ( .A1(p7_mult_21_n673), .A2(p7_mult_21_n691), .ZN(
        p7_mult_21_n379) );
  AOI21_X1 p7_mult_21_U492 ( .B1(p7_mult_21_n676), .B2(p7_mult_21_n674), .A(
        p7_mult_21_n690), .ZN(p7_mult_21_n689) );
  INV_X1 p7_mult_21_U491 ( .A(p7_mult_21_n689), .ZN(p7_mult_21_n380) );
  XNOR2_X1 p7_mult_21_U490 ( .A(B1[11]), .B(reg2_reg[5]), .ZN(p7_mult_21_n687)
         );
  OAI22_X1 p7_mult_21_U489 ( .A1(p7_mult_21_n687), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n688), .ZN(p7_mult_21_n381) );
  OAI22_X1 p7_mult_21_U488 ( .A1(p7_mult_21_n686), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n687), .ZN(p7_mult_21_n382) );
  XNOR2_X1 p7_mult_21_U487 ( .A(B1[8]), .B(reg2_reg[5]), .ZN(p7_mult_21_n684)
         );
  OAI22_X1 p7_mult_21_U486 ( .A1(p7_mult_21_n684), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n685), .ZN(p7_mult_21_n384) );
  XNOR2_X1 p7_mult_21_U485 ( .A(B1[7]), .B(reg2_reg[5]), .ZN(p7_mult_21_n683)
         );
  OAI22_X1 p7_mult_21_U484 ( .A1(p7_mult_21_n683), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n684), .ZN(p7_mult_21_n385) );
  XNOR2_X1 p7_mult_21_U483 ( .A(B1[6]), .B(reg2_reg[5]), .ZN(p7_mult_21_n682)
         );
  OAI22_X1 p7_mult_21_U482 ( .A1(p7_mult_21_n682), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n683), .ZN(p7_mult_21_n386) );
  XNOR2_X1 p7_mult_21_U481 ( .A(B1[5]), .B(reg2_reg[5]), .ZN(p7_mult_21_n681)
         );
  OAI22_X1 p7_mult_21_U480 ( .A1(p7_mult_21_n681), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n682), .ZN(p7_mult_21_n387) );
  XNOR2_X1 p7_mult_21_U479 ( .A(B1[4]), .B(reg2_reg[5]), .ZN(p7_mult_21_n680)
         );
  OAI22_X1 p7_mult_21_U478 ( .A1(p7_mult_21_n680), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n681), .ZN(p7_mult_21_n388) );
  XNOR2_X1 p7_mult_21_U477 ( .A(B1[3]), .B(reg2_reg[5]), .ZN(p7_mult_21_n679)
         );
  OAI22_X1 p7_mult_21_U476 ( .A1(p7_mult_21_n679), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n680), .ZN(p7_mult_21_n389) );
  XNOR2_X1 p7_mult_21_U475 ( .A(B1[2]), .B(reg2_reg[5]), .ZN(p7_mult_21_n678)
         );
  OAI22_X1 p7_mult_21_U474 ( .A1(p7_mult_21_n678), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n679), .ZN(p7_mult_21_n390) );
  XNOR2_X1 p7_mult_21_U473 ( .A(B1[1]), .B(reg2_reg[5]), .ZN(p7_mult_21_n677)
         );
  OAI22_X1 p7_mult_21_U472 ( .A1(p7_mult_21_n677), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n678), .ZN(p7_mult_21_n391) );
  XNOR2_X1 p7_mult_21_U471 ( .A(reg2_reg[5]), .B(B1[0]), .ZN(p7_mult_21_n675)
         );
  OAI22_X1 p7_mult_21_U470 ( .A1(p7_mult_21_n675), .A2(p7_mult_21_n676), .B1(
        p7_mult_21_n674), .B2(p7_mult_21_n677), .ZN(p7_mult_21_n392) );
  NOR2_X1 p7_mult_21_U469 ( .A1(p7_mult_21_n673), .A2(p7_mult_21_n674), .ZN(
        p7_mult_21_n393) );
  AOI21_X1 p7_mult_21_U468 ( .B1(p7_mult_21_n657), .B2(p7_mult_21_n658), .A(
        p7_mult_21_n672), .ZN(p7_mult_21_n671) );
  INV_X1 p7_mult_21_U467 ( .A(p7_mult_21_n671), .ZN(p7_mult_21_n394) );
  XNOR2_X1 p7_mult_21_U466 ( .A(B1[11]), .B(reg2_reg[3]), .ZN(p7_mult_21_n669)
         );
  OAI22_X1 p7_mult_21_U465 ( .A1(p7_mult_21_n669), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n670), .ZN(p7_mult_21_n395) );
  XNOR2_X1 p7_mult_21_U464 ( .A(B1[10]), .B(reg2_reg[3]), .ZN(p7_mult_21_n668)
         );
  OAI22_X1 p7_mult_21_U463 ( .A1(p7_mult_21_n668), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n669), .ZN(p7_mult_21_n396) );
  XNOR2_X1 p7_mult_21_U462 ( .A(B1[9]), .B(reg2_reg[3]), .ZN(p7_mult_21_n667)
         );
  OAI22_X1 p7_mult_21_U461 ( .A1(p7_mult_21_n667), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n668), .ZN(p7_mult_21_n397) );
  XNOR2_X1 p7_mult_21_U460 ( .A(B1[8]), .B(reg2_reg[3]), .ZN(p7_mult_21_n666)
         );
  OAI22_X1 p7_mult_21_U459 ( .A1(p7_mult_21_n666), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n667), .ZN(p7_mult_21_n398) );
  XNOR2_X1 p7_mult_21_U458 ( .A(B1[7]), .B(reg2_reg[3]), .ZN(p7_mult_21_n665)
         );
  OAI22_X1 p7_mult_21_U457 ( .A1(p7_mult_21_n665), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n666), .ZN(p7_mult_21_n399) );
  XNOR2_X1 p7_mult_21_U456 ( .A(B1[6]), .B(reg2_reg[3]), .ZN(p7_mult_21_n664)
         );
  OAI22_X1 p7_mult_21_U455 ( .A1(p7_mult_21_n664), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n665), .ZN(p7_mult_21_n400) );
  XNOR2_X1 p7_mult_21_U454 ( .A(B1[5]), .B(reg2_reg[3]), .ZN(p7_mult_21_n663)
         );
  OAI22_X1 p7_mult_21_U453 ( .A1(p7_mult_21_n663), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n664), .ZN(p7_mult_21_n401) );
  XNOR2_X1 p7_mult_21_U452 ( .A(B1[4]), .B(reg2_reg[3]), .ZN(p7_mult_21_n662)
         );
  OAI22_X1 p7_mult_21_U451 ( .A1(p7_mult_21_n662), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n663), .ZN(p7_mult_21_n402) );
  XNOR2_X1 p7_mult_21_U450 ( .A(B1[3]), .B(reg2_reg[3]), .ZN(p7_mult_21_n661)
         );
  OAI22_X1 p7_mult_21_U449 ( .A1(p7_mult_21_n661), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n662), .ZN(p7_mult_21_n403) );
  XNOR2_X1 p7_mult_21_U448 ( .A(B1[2]), .B(reg2_reg[3]), .ZN(p7_mult_21_n660)
         );
  OAI22_X1 p7_mult_21_U447 ( .A1(p7_mult_21_n660), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n661), .ZN(p7_mult_21_n404) );
  XNOR2_X1 p7_mult_21_U446 ( .A(B1[1]), .B(reg2_reg[3]), .ZN(p7_mult_21_n659)
         );
  OAI22_X1 p7_mult_21_U445 ( .A1(p7_mult_21_n659), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n660), .ZN(p7_mult_21_n405) );
  XNOR2_X1 p7_mult_21_U444 ( .A(reg2_reg[3]), .B(B1[0]), .ZN(p7_mult_21_n656)
         );
  OAI22_X1 p7_mult_21_U443 ( .A1(p7_mult_21_n656), .A2(p7_mult_21_n657), .B1(
        p7_mult_21_n658), .B2(p7_mult_21_n659), .ZN(p7_mult_21_n406) );
  XOR2_X1 p7_mult_21_U442 ( .A(B1[13]), .B(p7_mult_21_n655), .Z(
        p7_mult_21_n653) );
  AOI21_X1 p7_mult_21_U441 ( .B1(p7_mult_21_n641), .B2(p7_mult_21_n643), .A(
        p7_mult_21_n653), .ZN(p7_mult_21_n654) );
  INV_X1 p7_mult_21_U440 ( .A(p7_mult_21_n654), .ZN(p7_mult_21_n408) );
  XNOR2_X1 p7_mult_21_U439 ( .A(B1[12]), .B(reg2_reg[1]), .ZN(p7_mult_21_n652)
         );
  OAI22_X1 p7_mult_21_U438 ( .A1(p7_mult_21_n652), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n653), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n409) );
  XNOR2_X1 p7_mult_21_U437 ( .A(B1[11]), .B(reg2_reg[1]), .ZN(p7_mult_21_n651)
         );
  OAI22_X1 p7_mult_21_U436 ( .A1(p7_mult_21_n651), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n652), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n410) );
  XNOR2_X1 p7_mult_21_U435 ( .A(B1[10]), .B(reg2_reg[1]), .ZN(p7_mult_21_n650)
         );
  OAI22_X1 p7_mult_21_U434 ( .A1(p7_mult_21_n650), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n651), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n411) );
  XNOR2_X1 p7_mult_21_U433 ( .A(B1[9]), .B(reg2_reg[1]), .ZN(p7_mult_21_n649)
         );
  OAI22_X1 p7_mult_21_U432 ( .A1(p7_mult_21_n649), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n650), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n412) );
  XNOR2_X1 p7_mult_21_U431 ( .A(B1[8]), .B(reg2_reg[1]), .ZN(p7_mult_21_n648)
         );
  OAI22_X1 p7_mult_21_U430 ( .A1(p7_mult_21_n648), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n649), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n413) );
  XNOR2_X1 p7_mult_21_U429 ( .A(B1[7]), .B(reg2_reg[1]), .ZN(p7_mult_21_n647)
         );
  OAI22_X1 p7_mult_21_U428 ( .A1(p7_mult_21_n647), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n648), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n414) );
  XNOR2_X1 p7_mult_21_U427 ( .A(B1[6]), .B(reg2_reg[1]), .ZN(p7_mult_21_n646)
         );
  OAI22_X1 p7_mult_21_U426 ( .A1(p7_mult_21_n646), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n647), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n415) );
  XNOR2_X1 p7_mult_21_U425 ( .A(B1[5]), .B(reg2_reg[1]), .ZN(p7_mult_21_n645)
         );
  OAI22_X1 p7_mult_21_U424 ( .A1(p7_mult_21_n645), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n646), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n416) );
  XNOR2_X1 p7_mult_21_U423 ( .A(B1[4]), .B(reg2_reg[1]), .ZN(p7_mult_21_n644)
         );
  OAI22_X1 p7_mult_21_U422 ( .A1(p7_mult_21_n644), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n645), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n417) );
  XNOR2_X1 p7_mult_21_U421 ( .A(B1[3]), .B(reg2_reg[1]), .ZN(p7_mult_21_n642)
         );
  OAI22_X1 p7_mult_21_U420 ( .A1(p7_mult_21_n642), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n644), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n418) );
  OAI22_X1 p7_mult_21_U419 ( .A1(p7_mult_21_n640), .A2(p7_mult_21_n641), .B1(
        p7_mult_21_n642), .B2(p7_mult_21_n643), .ZN(p7_mult_21_n419) );
  OAI21_X1 p7_mult_21_U418 ( .B1(p7_mult_21_n637), .B2(p7_mult_21_n638), .A(
        p7_mult_21_n639), .ZN(p7_mult_21_n636) );
  XOR2_X1 p7_mult_21_U417 ( .A(p7_mult_21_n636), .B(p7_mult_21_n136), .Z(
        p7_mult_21_n635) );
  XNOR2_X1 p7_mult_21_U416 ( .A(p7_mult_21_n162), .B(p7_mult_21_n635), .ZN(
        temp2[13]) );
  XOR2_X2 p7_mult_21_U415 ( .A(reg2_reg[12]), .B(p7_mult_21_n764), .Z(
        p7_mult_21_n742) );
  XOR2_X2 p7_mult_21_U414 ( .A(reg2_reg[10]), .B(p7_mult_21_n762), .Z(
        p7_mult_21_n725) );
  XOR2_X2 p7_mult_21_U413 ( .A(reg2_reg[8]), .B(p7_mult_21_n760), .Z(
        p7_mult_21_n708) );
  XOR2_X2 p7_mult_21_U412 ( .A(reg2_reg[6]), .B(p7_mult_21_n758), .Z(
        p7_mult_21_n691) );
  XOR2_X2 p7_mult_21_U411 ( .A(reg2_reg[4]), .B(p7_mult_21_n771), .Z(
        p7_mult_21_n674) );
  INV_X1 p7_mult_21_U410 ( .A(reg2_reg[0]), .ZN(p7_mult_21_n643) );
  INV_X1 p7_mult_21_U409 ( .A(p7_mult_21_n798), .ZN(p7_mult_21_n658) );
  HA_X1 p7_mult_21_U145 ( .A(p7_mult_21_n406), .B(p7_mult_21_n419), .CO(
        p7_mult_21_n315), .S(p7_mult_21_n316) );
  FA_X1 p7_mult_21_U144 ( .A(p7_mult_21_n418), .B(p7_mult_21_n393), .CI(
        p7_mult_21_n405), .CO(p7_mult_21_n313), .S(p7_mult_21_n314) );
  HA_X1 p7_mult_21_U143 ( .A(p7_mult_21_n321), .B(p7_mult_21_n392), .CO(
        p7_mult_21_n311), .S(p7_mult_21_n312) );
  FA_X1 p7_mult_21_U142 ( .A(p7_mult_21_n404), .B(p7_mult_21_n417), .CI(
        p7_mult_21_n312), .CO(p7_mult_21_n309), .S(p7_mult_21_n310) );
  FA_X1 p7_mult_21_U141 ( .A(p7_mult_21_n416), .B(p7_mult_21_n379), .CI(
        p7_mult_21_n403), .CO(p7_mult_21_n307), .S(p7_mult_21_n308) );
  FA_X1 p7_mult_21_U140 ( .A(p7_mult_21_n311), .B(p7_mult_21_n391), .CI(
        p7_mult_21_n308), .CO(p7_mult_21_n305), .S(p7_mult_21_n306) );
  HA_X1 p7_mult_21_U139 ( .A(p7_mult_21_n320), .B(p7_mult_21_n378), .CO(
        p7_mult_21_n303), .S(p7_mult_21_n304) );
  FA_X1 p7_mult_21_U138 ( .A(p7_mult_21_n390), .B(p7_mult_21_n415), .CI(
        p7_mult_21_n402), .CO(p7_mult_21_n301), .S(p7_mult_21_n302) );
  FA_X1 p7_mult_21_U137 ( .A(p7_mult_21_n307), .B(p7_mult_21_n304), .CI(
        p7_mult_21_n302), .CO(p7_mult_21_n299), .S(p7_mult_21_n300) );
  FA_X1 p7_mult_21_U136 ( .A(p7_mult_21_n389), .B(p7_mult_21_n365), .CI(
        p7_mult_21_n414), .CO(p7_mult_21_n297), .S(p7_mult_21_n298) );
  FA_X1 p7_mult_21_U135 ( .A(p7_mult_21_n377), .B(p7_mult_21_n401), .CI(
        p7_mult_21_n303), .CO(p7_mult_21_n295), .S(p7_mult_21_n296) );
  FA_X1 p7_mult_21_U134 ( .A(p7_mult_21_n298), .B(p7_mult_21_n301), .CI(
        p7_mult_21_n296), .CO(p7_mult_21_n293), .S(p7_mult_21_n294) );
  HA_X1 p7_mult_21_U133 ( .A(p7_mult_21_n319), .B(p7_mult_21_n364), .CO(
        p7_mult_21_n291), .S(p7_mult_21_n292) );
  FA_X1 p7_mult_21_U132 ( .A(p7_mult_21_n376), .B(p7_mult_21_n388), .CI(
        p7_mult_21_n400), .CO(p7_mult_21_n289), .S(p7_mult_21_n290) );
  FA_X1 p7_mult_21_U131 ( .A(p7_mult_21_n292), .B(p7_mult_21_n413), .CI(
        p7_mult_21_n297), .CO(p7_mult_21_n287), .S(p7_mult_21_n288) );
  FA_X1 p7_mult_21_U130 ( .A(p7_mult_21_n290), .B(p7_mult_21_n295), .CI(
        p7_mult_21_n288), .CO(p7_mult_21_n285), .S(p7_mult_21_n286) );
  FA_X1 p7_mult_21_U129 ( .A(p7_mult_21_n375), .B(p7_mult_21_n351), .CI(
        p7_mult_21_n412), .CO(p7_mult_21_n283), .S(p7_mult_21_n284) );
  FA_X1 p7_mult_21_U128 ( .A(p7_mult_21_n363), .B(p7_mult_21_n399), .CI(
        p7_mult_21_n387), .CO(p7_mult_21_n281), .S(p7_mult_21_n282) );
  FA_X1 p7_mult_21_U127 ( .A(p7_mult_21_n289), .B(p7_mult_21_n291), .CI(
        p7_mult_21_n284), .CO(p7_mult_21_n279), .S(p7_mult_21_n280) );
  FA_X1 p7_mult_21_U126 ( .A(p7_mult_21_n287), .B(p7_mult_21_n282), .CI(
        p7_mult_21_n280), .CO(p7_mult_21_n277), .S(p7_mult_21_n278) );
  HA_X1 p7_mult_21_U125 ( .A(p7_mult_21_n318), .B(p7_mult_21_n350), .CO(
        p7_mult_21_n275), .S(p7_mult_21_n276) );
  FA_X1 p7_mult_21_U124 ( .A(p7_mult_21_n362), .B(p7_mult_21_n386), .CI(
        p7_mult_21_n411), .CO(p7_mult_21_n273), .S(p7_mult_21_n274) );
  FA_X1 p7_mult_21_U123 ( .A(p7_mult_21_n374), .B(p7_mult_21_n398), .CI(
        p7_mult_21_n276), .CO(p7_mult_21_n271), .S(p7_mult_21_n272) );
  FA_X1 p7_mult_21_U122 ( .A(p7_mult_21_n281), .B(p7_mult_21_n283), .CI(
        p7_mult_21_n274), .CO(p7_mult_21_n269), .S(p7_mult_21_n270) );
  FA_X1 p7_mult_21_U121 ( .A(p7_mult_21_n279), .B(p7_mult_21_n272), .CI(
        p7_mult_21_n270), .CO(p7_mult_21_n267), .S(p7_mult_21_n268) );
  FA_X1 p7_mult_21_U120 ( .A(p7_mult_21_n361), .B(p7_mult_21_n337), .CI(
        p7_mult_21_n410), .CO(p7_mult_21_n265), .S(p7_mult_21_n266) );
  FA_X1 p7_mult_21_U109 ( .A(p7_mult_21_n349), .B(p7_mult_21_n397), .CI(
        p7_mult_21_n373), .CO(p7_mult_21_n263), .S(p7_mult_21_n264) );
  FA_X1 p7_mult_21_U108 ( .A(p7_mult_21_n275), .B(p7_mult_21_n385), .CI(
        p7_mult_21_n273), .CO(p7_mult_21_n261), .S(p7_mult_21_n262) );
  FA_X1 p7_mult_21_U107 ( .A(p7_mult_21_n264), .B(p7_mult_21_n266), .CI(
        p7_mult_21_n271), .CO(p7_mult_21_n259), .S(p7_mult_21_n260) );
  FA_X1 p7_mult_21_U106 ( .A(p7_mult_21_n262), .B(p7_mult_21_n269), .CI(
        p7_mult_21_n260), .CO(p7_mult_21_n257), .S(p7_mult_21_n258) );
  HA_X1 p7_mult_21_U105 ( .A(p7_mult_21_n317), .B(p7_mult_21_n336), .CO(
        p7_mult_21_n255), .S(p7_mult_21_n256) );
  FA_X1 p7_mult_21_U104 ( .A(p7_mult_21_n409), .B(p7_mult_21_n372), .CI(
        p7_mult_21_n396), .CO(p7_mult_21_n253), .S(p7_mult_21_n254) );
  FA_X1 p7_mult_21_U103 ( .A(p7_mult_21_n348), .B(p7_mult_21_n384), .CI(
        p7_mult_21_n360), .CO(p7_mult_21_n251), .S(p7_mult_21_n252) );
  FA_X1 p7_mult_21_U102 ( .A(p7_mult_21_n265), .B(p7_mult_21_n256), .CI(
        p7_mult_21_n263), .CO(p7_mult_21_n249), .S(p7_mult_21_n250) );
  FA_X1 p7_mult_21_U101 ( .A(p7_mult_21_n254), .B(p7_mult_21_n252), .CI(
        p7_mult_21_n261), .CO(p7_mult_21_n247), .S(p7_mult_21_n248) );
  FA_X1 p7_mult_21_U100 ( .A(p7_mult_21_n259), .B(p7_mult_21_n250), .CI(
        p7_mult_21_n248), .CO(p7_mult_21_n245), .S(p7_mult_21_n246) );
  FA_X1 p7_mult_21_U97 ( .A(p7_mult_21_n395), .B(p7_mult_21_n359), .CI(
        p7_mult_21_n408), .CO(p7_mult_21_n241), .S(p7_mult_21_n242) );
  FA_X1 p7_mult_21_U96 ( .A(p7_mult_21_n335), .B(p7_mult_21_n371), .CI(
        p7_mult_21_n255), .CO(p7_mult_21_n239), .S(p7_mult_21_n240) );
  FA_X1 p7_mult_21_U95 ( .A(p7_mult_21_n253), .B(p7_mult_21_n244), .CI(
        p7_mult_21_n251), .CO(p7_mult_21_n237), .S(p7_mult_21_n238) );
  FA_X1 p7_mult_21_U94 ( .A(p7_mult_21_n240), .B(p7_mult_21_n242), .CI(
        p7_mult_21_n249), .CO(p7_mult_21_n235), .S(p7_mult_21_n236) );
  FA_X1 p7_mult_21_U93 ( .A(p7_mult_21_n247), .B(p7_mult_21_n238), .CI(
        p7_mult_21_n236), .CO(p7_mult_21_n233), .S(p7_mult_21_n234) );
  FA_X1 p7_mult_21_U91 ( .A(p7_mult_21_n382), .B(p7_mult_21_n346), .CI(
        p7_mult_21_n232), .CO(p7_mult_21_n229), .S(p7_mult_21_n230) );
  FA_X1 p7_mult_21_U90 ( .A(p7_mult_21_n334), .B(p7_mult_21_n370), .CI(
        p7_mult_21_n358), .CO(p7_mult_21_n227), .S(p7_mult_21_n228) );
  FA_X1 p7_mult_21_U89 ( .A(p7_mult_21_n241), .B(p7_mult_21_n243), .CI(
        p7_mult_21_n239), .CO(p7_mult_21_n225), .S(p7_mult_21_n226) );
  FA_X1 p7_mult_21_U88 ( .A(p7_mult_21_n230), .B(p7_mult_21_n228), .CI(
        p7_mult_21_n237), .CO(p7_mult_21_n223), .S(p7_mult_21_n224) );
  FA_X1 p7_mult_21_U87 ( .A(p7_mult_21_n235), .B(p7_mult_21_n226), .CI(
        p7_mult_21_n224), .CO(p7_mult_21_n221), .S(p7_mult_21_n222) );
  FA_X1 p7_mult_21_U86 ( .A(p7_mult_21_n231), .B(p7_mult_21_n333), .CI(
        p7_mult_21_n394), .CO(p7_mult_21_n219), .S(p7_mult_21_n220) );
  FA_X1 p7_mult_21_U85 ( .A(p7_mult_21_n345), .B(p7_mult_21_n381), .CI(
        p7_mult_21_n357), .CO(p7_mult_21_n217), .S(p7_mult_21_n218) );
  FA_X1 p7_mult_21_U84 ( .A(p7_mult_21_n229), .B(p7_mult_21_n369), .CI(
        p7_mult_21_n227), .CO(p7_mult_21_n215), .S(p7_mult_21_n216) );
  FA_X1 p7_mult_21_U83 ( .A(p7_mult_21_n220), .B(p7_mult_21_n218), .CI(
        p7_mult_21_n225), .CO(p7_mult_21_n213), .S(p7_mult_21_n214) );
  FA_X1 p7_mult_21_U82 ( .A(p7_mult_21_n223), .B(p7_mult_21_n216), .CI(
        p7_mult_21_n214), .CO(p7_mult_21_n211), .S(p7_mult_21_n212) );
  FA_X1 p7_mult_21_U80 ( .A(p7_mult_21_n368), .B(p7_mult_21_n344), .CI(
        p7_mult_21_n210), .CO(p7_mult_21_n207), .S(p7_mult_21_n208) );
  FA_X1 p7_mult_21_U79 ( .A(p7_mult_21_n332), .B(p7_mult_21_n356), .CI(
        p7_mult_21_n219), .CO(p7_mult_21_n205), .S(p7_mult_21_n206) );
  FA_X1 p7_mult_21_U78 ( .A(p7_mult_21_n208), .B(p7_mult_21_n217), .CI(
        p7_mult_21_n215), .CO(p7_mult_21_n203), .S(p7_mult_21_n204) );
  FA_X1 p7_mult_21_U77 ( .A(p7_mult_21_n213), .B(p7_mult_21_n206), .CI(
        p7_mult_21_n204), .CO(p7_mult_21_n201), .S(p7_mult_21_n202) );
  FA_X1 p7_mult_21_U76 ( .A(p7_mult_21_n209), .B(p7_mult_21_n331), .CI(
        p7_mult_21_n380), .CO(p7_mult_21_n199), .S(p7_mult_21_n200) );
  FA_X1 p7_mult_21_U75 ( .A(p7_mult_21_n355), .B(p7_mult_21_n343), .CI(
        p7_mult_21_n367), .CO(p7_mult_21_n197), .S(p7_mult_21_n198) );
  FA_X1 p7_mult_21_U74 ( .A(p7_mult_21_n198), .B(p7_mult_21_n207), .CI(
        p7_mult_21_n200), .CO(p7_mult_21_n195), .S(p7_mult_21_n196) );
  FA_X1 p7_mult_21_U73 ( .A(p7_mult_21_n203), .B(p7_mult_21_n205), .CI(
        p7_mult_21_n196), .CO(p7_mult_21_n193), .S(p7_mult_21_n194) );
  FA_X1 p7_mult_21_U71 ( .A(p7_mult_21_n330), .B(p7_mult_21_n342), .CI(
        p7_mult_21_n192), .CO(p7_mult_21_n189), .S(p7_mult_21_n190) );
  FA_X1 p7_mult_21_U70 ( .A(p7_mult_21_n199), .B(p7_mult_21_n354), .CI(
        p7_mult_21_n197), .CO(p7_mult_21_n187), .S(p7_mult_21_n188) );
  FA_X1 p7_mult_21_U69 ( .A(p7_mult_21_n188), .B(p7_mult_21_n190), .CI(
        p7_mult_21_n195), .CO(p7_mult_21_n185), .S(p7_mult_21_n186) );
  FA_X1 p7_mult_21_U68 ( .A(p7_mult_21_n191), .B(p7_mult_21_n329), .CI(
        p7_mult_21_n366), .CO(p7_mult_21_n183), .S(p7_mult_21_n184) );
  FA_X1 p7_mult_21_U67 ( .A(p7_mult_21_n341), .B(p7_mult_21_n353), .CI(
        p7_mult_21_n189), .CO(p7_mult_21_n181), .S(p7_mult_21_n182) );
  FA_X1 p7_mult_21_U66 ( .A(p7_mult_21_n187), .B(p7_mult_21_n184), .CI(
        p7_mult_21_n182), .CO(p7_mult_21_n179), .S(p7_mult_21_n180) );
  FA_X1 p7_mult_21_U64 ( .A(p7_mult_21_n328), .B(p7_mult_21_n340), .CI(
        p7_mult_21_n178), .CO(p7_mult_21_n175), .S(p7_mult_21_n176) );
  FA_X1 p7_mult_21_U63 ( .A(p7_mult_21_n176), .B(p7_mult_21_n183), .CI(
        p7_mult_21_n181), .CO(p7_mult_21_n173), .S(p7_mult_21_n174) );
  FA_X1 p7_mult_21_U62 ( .A(p7_mult_21_n327), .B(p7_mult_21_n177), .CI(
        p7_mult_21_n352), .CO(p7_mult_21_n171), .S(p7_mult_21_n172) );
  FA_X1 p7_mult_21_U61 ( .A(p7_mult_21_n175), .B(p7_mult_21_n339), .CI(
        p7_mult_21_n172), .CO(p7_mult_21_n169), .S(p7_mult_21_n170) );
  FA_X1 p7_mult_21_U59 ( .A(p7_mult_21_n168), .B(p7_mult_21_n326), .CI(
        p7_mult_21_n171), .CO(p7_mult_21_n165), .S(p7_mult_21_n166) );
  FA_X1 p7_mult_21_U58 ( .A(p7_mult_21_n325), .B(p7_mult_21_n167), .CI(
        p7_mult_21_n338), .CO(p7_mult_21_n163), .S(p7_mult_21_n164) );
  FA_X1 p7_mult_21_U44 ( .A(p7_mult_21_n246), .B(p7_mult_21_n257), .CI(
        p7_mult_21_n149), .CO(p7_mult_21_n148), .S(temp2[0]) );
  FA_X1 p7_mult_21_U43 ( .A(p7_mult_21_n234), .B(p7_mult_21_n245), .CI(
        p7_mult_21_n148), .CO(p7_mult_21_n147), .S(temp2[1]) );
  FA_X1 p7_mult_21_U42 ( .A(p7_mult_21_n222), .B(p7_mult_21_n233), .CI(
        p7_mult_21_n147), .CO(p7_mult_21_n146), .S(temp2[2]) );
  FA_X1 p7_mult_21_U41 ( .A(p7_mult_21_n212), .B(p7_mult_21_n221), .CI(
        p7_mult_21_n146), .CO(p7_mult_21_n145), .S(temp2[3]) );
  FA_X1 p7_mult_21_U40 ( .A(p7_mult_21_n202), .B(p7_mult_21_n211), .CI(
        p7_mult_21_n145), .CO(p7_mult_21_n144), .S(temp2[4]) );
  FA_X1 p7_mult_21_U39 ( .A(p7_mult_21_n194), .B(p7_mult_21_n201), .CI(
        p7_mult_21_n144), .CO(p7_mult_21_n143), .S(temp2[5]) );
  FA_X1 p7_mult_21_U38 ( .A(p7_mult_21_n186), .B(p7_mult_21_n193), .CI(
        p7_mult_21_n143), .CO(p7_mult_21_n142), .S(temp2[6]) );
  FA_X1 p7_mult_21_U37 ( .A(p7_mult_21_n180), .B(p7_mult_21_n185), .CI(
        p7_mult_21_n142), .CO(p7_mult_21_n141), .S(temp2[7]) );
  FA_X1 p7_mult_21_U30 ( .A(p7_mult_21_n174), .B(p7_mult_21_n179), .CI(
        p7_mult_21_n141), .CO(p7_mult_21_n140), .S(temp2[8]) );
  FA_X1 p7_mult_21_U20 ( .A(p7_mult_21_n170), .B(p7_mult_21_n173), .CI(
        p7_mult_21_n140), .CO(p7_mult_21_n139), .S(temp2[9]) );
  FA_X1 p7_mult_21_U10 ( .A(p7_mult_21_n166), .B(p7_mult_21_n169), .CI(
        p7_mult_21_n139), .CO(p7_mult_21_n138), .S(temp2[10]) );
  FA_X1 p7_mult_21_U9 ( .A(p7_mult_21_n165), .B(p7_mult_21_n164), .CI(
        p7_mult_21_n138), .CO(p7_mult_21_n137), .S(temp2[11]) );
  FA_X1 p7_mult_21_U8 ( .A(p7_mult_21_n163), .B(p7_mult_21_n162), .CI(
        p7_mult_21_n137), .CO(p7_mult_21_n136), .S(temp2[12]) );
  NAND2_X1 REG2_1_U34 ( .A1(temp2[4]), .A2(REG2_1_n43), .ZN(REG2_1_n85) );
  OAI21_X1 REG2_1_U33 ( .B1(REG2_1_n45), .B2(REG2_1_n66), .A(REG2_1_n85), .ZN(
        REG2_1_n57) );
  NAND2_X1 REG2_1_U32 ( .A1(temp2[3]), .A2(REG2_1_n43), .ZN(REG2_1_n86) );
  OAI21_X1 REG2_1_U31 ( .B1(REG2_1_n45), .B2(REG2_1_n65), .A(REG2_1_n86), .ZN(
        REG2_1_n58) );
  NAND2_X1 REG2_1_U30 ( .A1(temp2[2]), .A2(REG2_1_n43), .ZN(REG2_1_n87) );
  OAI21_X1 REG2_1_U29 ( .B1(REG2_1_n45), .B2(REG2_1_n64), .A(REG2_1_n87), .ZN(
        REG2_1_n59) );
  NAND2_X1 REG2_1_U28 ( .A1(temp2[5]), .A2(REG2_1_n43), .ZN(REG2_1_n84) );
  OAI21_X1 REG2_1_U27 ( .B1(REG2_1_n44), .B2(REG2_1_n67), .A(REG2_1_n84), .ZN(
        REG2_1_n56) );
  NAND2_X1 REG2_1_U26 ( .A1(temp2[9]), .A2(REG2_1_n43), .ZN(REG2_1_n80) );
  OAI21_X1 REG2_1_U25 ( .B1(REG2_1_n44), .B2(REG2_1_n71), .A(REG2_1_n80), .ZN(
        REG2_1_n52) );
  NAND2_X1 REG2_1_U24 ( .A1(temp2[8]), .A2(REG2_1_n44), .ZN(REG2_1_n81) );
  OAI21_X1 REG2_1_U23 ( .B1(REG2_1_n44), .B2(REG2_1_n70), .A(REG2_1_n81), .ZN(
        REG2_1_n53) );
  NAND2_X1 REG2_1_U22 ( .A1(temp2[7]), .A2(REG2_1_n43), .ZN(REG2_1_n82) );
  OAI21_X1 REG2_1_U21 ( .B1(REG2_1_n44), .B2(REG2_1_n69), .A(REG2_1_n82), .ZN(
        REG2_1_n54) );
  NAND2_X1 REG2_1_U20 ( .A1(temp2[6]), .A2(REG2_1_n43), .ZN(REG2_1_n83) );
  OAI21_X1 REG2_1_U19 ( .B1(REG2_1_n44), .B2(REG2_1_n68), .A(REG2_1_n83), .ZN(
        REG2_1_n55) );
  NAND2_X1 REG2_1_U18 ( .A1(temp2[1]), .A2(REG2_1_n43), .ZN(REG2_1_n88) );
  OAI21_X1 REG2_1_U17 ( .B1(REG2_1_n44), .B2(REG2_1_n63), .A(REG2_1_n88), .ZN(
        REG2_1_n60) );
  NAND2_X1 REG2_1_U16 ( .A1(temp2[0]), .A2(REG2_1_n43), .ZN(REG2_1_n89) );
  OAI21_X1 REG2_1_U15 ( .B1(REG2_1_n44), .B2(REG2_1_n62), .A(REG2_1_n89), .ZN(
        REG2_1_n61) );
  NAND2_X1 REG2_1_U14 ( .A1(temp2[10]), .A2(REG2_1_n44), .ZN(REG2_1_n79) );
  OAI21_X1 REG2_1_U13 ( .B1(REG2_1_n44), .B2(REG2_1_n72), .A(REG2_1_n79), .ZN(
        REG2_1_n51) );
  NAND2_X1 REG2_1_U12 ( .A1(temp2[12]), .A2(REG2_1_n43), .ZN(REG2_1_n77) );
  OAI21_X1 REG2_1_U11 ( .B1(REG2_1_n44), .B2(REG2_1_n74), .A(REG2_1_n77), .ZN(
        REG2_1_n49) );
  NAND2_X1 REG2_1_U10 ( .A1(temp2[11]), .A2(REG2_1_n43), .ZN(REG2_1_n78) );
  OAI21_X1 REG2_1_U9 ( .B1(REG2_1_n44), .B2(REG2_1_n73), .A(REG2_1_n78), .ZN(
        REG2_1_n50) );
  NAND2_X1 REG2_1_U8 ( .A1(temp2[13]), .A2(REG2_1_n43), .ZN(REG2_1_n76) );
  OAI21_X1 REG2_1_U7 ( .B1(REG2_1_n44), .B2(REG2_1_n75), .A(REG2_1_n76), .ZN(
        REG2_1_n48) );
  BUF_X1 REG2_1_U6 ( .A(n47), .Z(REG2_1_n47) );
  BUF_X1 REG2_1_U5 ( .A(n47), .Z(REG2_1_n46) );
  BUF_X1 REG2_1_U4 ( .A(VIN), .Z(REG2_1_n45) );
  BUF_X1 REG2_1_U3 ( .A(VIN), .Z(REG2_1_n43) );
  BUF_X1 REG2_1_U2 ( .A(VIN), .Z(REG2_1_n44) );
  DFFR_X1 REG2_1_q_reg_0_ ( .D(REG2_1_n61), .CK(CLK), .RN(REG2_1_n47), .Q(
        mul2_reg[0]), .QN(REG2_1_n62) );
  DFFR_X1 REG2_1_q_reg_1_ ( .D(REG2_1_n60), .CK(CLK), .RN(REG2_1_n47), .Q(
        mul2_reg[1]), .QN(REG2_1_n63) );
  DFFR_X1 REG2_1_q_reg_2_ ( .D(REG2_1_n59), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[2]), .QN(REG2_1_n64) );
  DFFR_X1 REG2_1_q_reg_3_ ( .D(REG2_1_n58), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[3]), .QN(REG2_1_n65) );
  DFFR_X1 REG2_1_q_reg_4_ ( .D(REG2_1_n57), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[4]), .QN(REG2_1_n66) );
  DFFR_X1 REG2_1_q_reg_5_ ( .D(REG2_1_n56), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[5]), .QN(REG2_1_n67) );
  DFFR_X1 REG2_1_q_reg_6_ ( .D(REG2_1_n55), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[6]), .QN(REG2_1_n68) );
  DFFR_X1 REG2_1_q_reg_7_ ( .D(REG2_1_n54), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[7]), .QN(REG2_1_n69) );
  DFFR_X1 REG2_1_q_reg_8_ ( .D(REG2_1_n53), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[8]), .QN(REG2_1_n70) );
  DFFR_X1 REG2_1_q_reg_9_ ( .D(REG2_1_n52), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[9]), .QN(REG2_1_n71) );
  DFFR_X1 REG2_1_q_reg_10_ ( .D(REG2_1_n51), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[10]), .QN(REG2_1_n72) );
  DFFR_X1 REG2_1_q_reg_11_ ( .D(REG2_1_n50), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[11]), .QN(REG2_1_n73) );
  DFFR_X1 REG2_1_q_reg_12_ ( .D(REG2_1_n49), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[12]), .QN(REG2_1_n74) );
  DFFR_X1 REG2_1_q_reg_13_ ( .D(REG2_1_n48), .CK(CLK), .RN(REG2_1_n46), .Q(
        mul2_reg[13]), .QN(REG2_1_n75) );
  NAND2_X1 REGISTER3_U34 ( .A1(reg3[13]), .A2(REGISTER3_n43), .ZN(
        REGISTER3_n76) );
  OAI21_X1 REGISTER3_U33 ( .B1(REGISTER3_n44), .B2(REGISTER3_n75), .A(
        REGISTER3_n76), .ZN(REGISTER3_n48) );
  NAND2_X1 REGISTER3_U32 ( .A1(reg3[12]), .A2(REGISTER3_n43), .ZN(
        REGISTER3_n77) );
  OAI21_X1 REGISTER3_U31 ( .B1(REGISTER3_n44), .B2(REGISTER3_n74), .A(
        REGISTER3_n77), .ZN(REGISTER3_n49) );
  NAND2_X1 REGISTER3_U30 ( .A1(reg3[11]), .A2(REGISTER3_n43), .ZN(
        REGISTER3_n78) );
  OAI21_X1 REGISTER3_U29 ( .B1(REGISTER3_n44), .B2(REGISTER3_n73), .A(
        REGISTER3_n78), .ZN(REGISTER3_n50) );
  NAND2_X1 REGISTER3_U28 ( .A1(reg3[9]), .A2(REGISTER3_n43), .ZN(REGISTER3_n80) );
  OAI21_X1 REGISTER3_U27 ( .B1(REGISTER3_n44), .B2(REGISTER3_n71), .A(
        REGISTER3_n80), .ZN(REGISTER3_n52) );
  NAND2_X1 REGISTER3_U26 ( .A1(reg3[7]), .A2(REGISTER3_n43), .ZN(REGISTER3_n82) );
  OAI21_X1 REGISTER3_U25 ( .B1(REGISTER3_n44), .B2(REGISTER3_n69), .A(
        REGISTER3_n82), .ZN(REGISTER3_n54) );
  NAND2_X1 REGISTER3_U24 ( .A1(reg3[6]), .A2(REGISTER3_n43), .ZN(REGISTER3_n83) );
  OAI21_X1 REGISTER3_U23 ( .B1(REGISTER3_n44), .B2(REGISTER3_n68), .A(
        REGISTER3_n83), .ZN(REGISTER3_n55) );
  NAND2_X1 REGISTER3_U22 ( .A1(reg3[5]), .A2(REGISTER3_n43), .ZN(REGISTER3_n84) );
  OAI21_X1 REGISTER3_U21 ( .B1(REGISTER3_n44), .B2(REGISTER3_n67), .A(
        REGISTER3_n84), .ZN(REGISTER3_n56) );
  NAND2_X1 REGISTER3_U20 ( .A1(reg3[4]), .A2(REGISTER3_n43), .ZN(REGISTER3_n85) );
  OAI21_X1 REGISTER3_U19 ( .B1(REGISTER3_n45), .B2(REGISTER3_n66), .A(
        REGISTER3_n85), .ZN(REGISTER3_n57) );
  NAND2_X1 REGISTER3_U18 ( .A1(reg3[3]), .A2(REGISTER3_n43), .ZN(REGISTER3_n86) );
  OAI21_X1 REGISTER3_U17 ( .B1(REGISTER3_n45), .B2(REGISTER3_n65), .A(
        REGISTER3_n86), .ZN(REGISTER3_n58) );
  NAND2_X1 REGISTER3_U16 ( .A1(reg3[2]), .A2(REGISTER3_n43), .ZN(REGISTER3_n87) );
  OAI21_X1 REGISTER3_U15 ( .B1(REGISTER3_n45), .B2(REGISTER3_n64), .A(
        REGISTER3_n87), .ZN(REGISTER3_n59) );
  NAND2_X1 REGISTER3_U14 ( .A1(reg3[1]), .A2(REGISTER3_n43), .ZN(REGISTER3_n88) );
  OAI21_X1 REGISTER3_U13 ( .B1(REGISTER3_n44), .B2(REGISTER3_n63), .A(
        REGISTER3_n88), .ZN(REGISTER3_n60) );
  NAND2_X1 REGISTER3_U12 ( .A1(reg3[0]), .A2(REGISTER3_n43), .ZN(REGISTER3_n89) );
  OAI21_X1 REGISTER3_U11 ( .B1(REGISTER3_n44), .B2(REGISTER3_n62), .A(
        REGISTER3_n89), .ZN(REGISTER3_n61) );
  NAND2_X1 REGISTER3_U10 ( .A1(reg3[10]), .A2(REGISTER3_n44), .ZN(
        REGISTER3_n79) );
  OAI21_X1 REGISTER3_U9 ( .B1(REGISTER3_n44), .B2(REGISTER3_n72), .A(
        REGISTER3_n79), .ZN(REGISTER3_n51) );
  NAND2_X1 REGISTER3_U8 ( .A1(reg3[8]), .A2(REGISTER3_n44), .ZN(REGISTER3_n81)
         );
  OAI21_X1 REGISTER3_U7 ( .B1(REGISTER3_n44), .B2(REGISTER3_n70), .A(
        REGISTER3_n81), .ZN(REGISTER3_n53) );
  BUF_X1 REGISTER3_U6 ( .A(n47), .Z(REGISTER3_n47) );
  BUF_X1 REGISTER3_U5 ( .A(n47), .Z(REGISTER3_n46) );
  BUF_X1 REGISTER3_U4 ( .A(VIN), .Z(REGISTER3_n45) );
  BUF_X1 REGISTER3_U3 ( .A(VIN), .Z(REGISTER3_n43) );
  BUF_X1 REGISTER3_U2 ( .A(VIN), .Z(REGISTER3_n44) );
  DFFR_X1 REGISTER3_q_reg_0_ ( .D(REGISTER3_n61), .CK(CLK), .RN(REGISTER3_n47), 
        .Q(reg3_reg[0]), .QN(REGISTER3_n62) );
  DFFR_X1 REGISTER3_q_reg_1_ ( .D(REGISTER3_n60), .CK(CLK), .RN(REGISTER3_n47), 
        .Q(reg3_reg[1]), .QN(REGISTER3_n63) );
  DFFR_X1 REGISTER3_q_reg_2_ ( .D(REGISTER3_n59), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[2]), .QN(REGISTER3_n64) );
  DFFR_X1 REGISTER3_q_reg_3_ ( .D(REGISTER3_n58), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[3]), .QN(REGISTER3_n65) );
  DFFR_X1 REGISTER3_q_reg_4_ ( .D(REGISTER3_n57), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[4]), .QN(REGISTER3_n66) );
  DFFR_X1 REGISTER3_q_reg_5_ ( .D(REGISTER3_n56), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[5]), .QN(REGISTER3_n67) );
  DFFR_X1 REGISTER3_q_reg_6_ ( .D(REGISTER3_n55), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[6]), .QN(REGISTER3_n68) );
  DFFR_X1 REGISTER3_q_reg_7_ ( .D(REGISTER3_n54), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[7]), .QN(REGISTER3_n69) );
  DFFR_X1 REGISTER3_q_reg_8_ ( .D(REGISTER3_n53), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[8]), .QN(REGISTER3_n70) );
  DFFR_X1 REGISTER3_q_reg_9_ ( .D(REGISTER3_n52), .CK(CLK), .RN(REGISTER3_n46), 
        .Q(reg3_reg[9]), .QN(REGISTER3_n71) );
  DFFR_X1 REGISTER3_q_reg_10_ ( .D(REGISTER3_n51), .CK(CLK), .RN(REGISTER3_n46), .Q(reg3_reg[10]), .QN(REGISTER3_n72) );
  DFFR_X1 REGISTER3_q_reg_11_ ( .D(REGISTER3_n50), .CK(CLK), .RN(REGISTER3_n46), .Q(reg3_reg[11]), .QN(REGISTER3_n73) );
  DFFR_X1 REGISTER3_q_reg_12_ ( .D(REGISTER3_n49), .CK(CLK), .RN(REGISTER3_n46), .Q(reg3_reg[12]), .QN(REGISTER3_n74) );
  DFFR_X1 REGISTER3_q_reg_13_ ( .D(REGISTER3_n48), .CK(CLK), .RN(REGISTER3_n46), .Q(reg3_reg[13]), .QN(REGISTER3_n75) );
  XOR2_X1 p8_mult_21_U691 ( .A(reg3_reg[2]), .B(reg3_reg[1]), .Z(
        p8_mult_21_n798) );
  INV_X1 p8_mult_21_U690 ( .A(reg3_reg[1]), .ZN(p8_mult_21_n655) );
  NOR2_X1 p8_mult_21_U689 ( .A1(p8_mult_21_n655), .A2(B2[1]), .ZN(
        p8_mult_21_n803) );
  INV_X1 p8_mult_21_U688 ( .A(p8_mult_21_n803), .ZN(p8_mult_21_n805) );
  NAND2_X1 p8_mult_21_U687 ( .A1(reg3_reg[1]), .A2(p8_mult_21_n643), .ZN(
        p8_mult_21_n641) );
  XNOR2_X1 p8_mult_21_U686 ( .A(B2[2]), .B(reg3_reg[1]), .ZN(p8_mult_21_n640)
         );
  OAI22_X1 p8_mult_21_U685 ( .A1(p8_mult_21_n805), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n640), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n804) );
  NAND2_X1 p8_mult_21_U684 ( .A1(p8_mult_21_n798), .A2(p8_mult_21_n804), .ZN(
        p8_mult_21_n801) );
  NAND2_X1 p8_mult_21_U683 ( .A1(p8_mult_21_n803), .A2(p8_mult_21_n804), .ZN(
        p8_mult_21_n802) );
  INV_X1 p8_mult_21_U682 ( .A(B2[0]), .ZN(p8_mult_21_n673) );
  MUX2_X1 p8_mult_21_U681 ( .A(p8_mult_21_n801), .B(p8_mult_21_n802), .S(
        p8_mult_21_n673), .Z(p8_mult_21_n800) );
  INV_X1 p8_mult_21_U680 ( .A(p8_mult_21_n800), .ZN(p8_mult_21_n795) );
  INV_X1 p8_mult_21_U679 ( .A(reg3_reg[3]), .ZN(p8_mult_21_n771) );
  XNOR2_X1 p8_mult_21_U678 ( .A(p8_mult_21_n771), .B(reg3_reg[2]), .ZN(
        p8_mult_21_n799) );
  NAND2_X1 p8_mult_21_U677 ( .A1(p8_mult_21_n658), .A2(p8_mult_21_n799), .ZN(
        p8_mult_21_n657) );
  NAND3_X1 p8_mult_21_U676 ( .A1(p8_mult_21_n798), .A2(p8_mult_21_n673), .A3(
        reg3_reg[3]), .ZN(p8_mult_21_n797) );
  OAI21_X1 p8_mult_21_U675 ( .B1(p8_mult_21_n771), .B2(p8_mult_21_n657), .A(
        p8_mult_21_n797), .ZN(p8_mult_21_n796) );
  AOI222_X1 p8_mult_21_U674 ( .A1(p8_mult_21_n795), .A2(p8_mult_21_n316), .B1(
        p8_mult_21_n796), .B2(p8_mult_21_n795), .C1(p8_mult_21_n796), .C2(
        p8_mult_21_n316), .ZN(p8_mult_21_n794) );
  INV_X1 p8_mult_21_U673 ( .A(p8_mult_21_n794), .ZN(p8_mult_21_n793) );
  AOI222_X1 p8_mult_21_U672 ( .A1(p8_mult_21_n793), .A2(p8_mult_21_n314), .B1(
        p8_mult_21_n793), .B2(p8_mult_21_n315), .C1(p8_mult_21_n315), .C2(
        p8_mult_21_n314), .ZN(p8_mult_21_n792) );
  INV_X1 p8_mult_21_U671 ( .A(p8_mult_21_n792), .ZN(p8_mult_21_n791) );
  AOI222_X1 p8_mult_21_U670 ( .A1(p8_mult_21_n791), .A2(p8_mult_21_n310), .B1(
        p8_mult_21_n791), .B2(p8_mult_21_n313), .C1(p8_mult_21_n313), .C2(
        p8_mult_21_n310), .ZN(p8_mult_21_n790) );
  INV_X1 p8_mult_21_U669 ( .A(p8_mult_21_n790), .ZN(p8_mult_21_n789) );
  AOI222_X1 p8_mult_21_U668 ( .A1(p8_mult_21_n789), .A2(p8_mult_21_n306), .B1(
        p8_mult_21_n789), .B2(p8_mult_21_n309), .C1(p8_mult_21_n309), .C2(
        p8_mult_21_n306), .ZN(p8_mult_21_n788) );
  INV_X1 p8_mult_21_U667 ( .A(p8_mult_21_n788), .ZN(p8_mult_21_n787) );
  AOI222_X1 p8_mult_21_U666 ( .A1(p8_mult_21_n787), .A2(p8_mult_21_n300), .B1(
        p8_mult_21_n787), .B2(p8_mult_21_n305), .C1(p8_mult_21_n305), .C2(
        p8_mult_21_n300), .ZN(p8_mult_21_n786) );
  INV_X1 p8_mult_21_U665 ( .A(p8_mult_21_n786), .ZN(p8_mult_21_n785) );
  AOI222_X1 p8_mult_21_U664 ( .A1(p8_mult_21_n785), .A2(p8_mult_21_n294), .B1(
        p8_mult_21_n785), .B2(p8_mult_21_n299), .C1(p8_mult_21_n299), .C2(
        p8_mult_21_n294), .ZN(p8_mult_21_n784) );
  INV_X1 p8_mult_21_U663 ( .A(p8_mult_21_n784), .ZN(p8_mult_21_n783) );
  AOI222_X1 p8_mult_21_U662 ( .A1(p8_mult_21_n783), .A2(p8_mult_21_n286), .B1(
        p8_mult_21_n783), .B2(p8_mult_21_n293), .C1(p8_mult_21_n293), .C2(
        p8_mult_21_n286), .ZN(p8_mult_21_n780) );
  INV_X1 p8_mult_21_U661 ( .A(p8_mult_21_n278), .ZN(p8_mult_21_n781) );
  INV_X1 p8_mult_21_U660 ( .A(p8_mult_21_n285), .ZN(p8_mult_21_n782) );
  OAI222_X1 p8_mult_21_U659 ( .A1(p8_mult_21_n780), .A2(p8_mult_21_n781), .B1(
        p8_mult_21_n780), .B2(p8_mult_21_n782), .C1(p8_mult_21_n782), .C2(
        p8_mult_21_n781), .ZN(p8_mult_21_n779) );
  AOI222_X1 p8_mult_21_U658 ( .A1(p8_mult_21_n779), .A2(p8_mult_21_n268), .B1(
        p8_mult_21_n779), .B2(p8_mult_21_n277), .C1(p8_mult_21_n277), .C2(
        p8_mult_21_n268), .ZN(p8_mult_21_n776) );
  INV_X1 p8_mult_21_U657 ( .A(p8_mult_21_n258), .ZN(p8_mult_21_n777) );
  INV_X1 p8_mult_21_U656 ( .A(p8_mult_21_n267), .ZN(p8_mult_21_n778) );
  OAI222_X1 p8_mult_21_U655 ( .A1(p8_mult_21_n776), .A2(p8_mult_21_n777), .B1(
        p8_mult_21_n776), .B2(p8_mult_21_n778), .C1(p8_mult_21_n778), .C2(
        p8_mult_21_n777), .ZN(p8_mult_21_n149) );
  XOR2_X1 p8_mult_21_U654 ( .A(B2[12]), .B(reg3_reg[13]), .Z(p8_mult_21_n757)
         );
  INV_X1 p8_mult_21_U653 ( .A(reg3_reg[11]), .ZN(p8_mult_21_n764) );
  INV_X1 p8_mult_21_U652 ( .A(reg3_reg[13]), .ZN(p8_mult_21_n766) );
  XNOR2_X1 p8_mult_21_U651 ( .A(p8_mult_21_n766), .B(reg3_reg[12]), .ZN(
        p8_mult_21_n775) );
  NAND2_X1 p8_mult_21_U650 ( .A1(p8_mult_21_n742), .A2(p8_mult_21_n775), .ZN(
        p8_mult_21_n744) );
  INV_X1 p8_mult_21_U649 ( .A(p8_mult_21_n744), .ZN(p8_mult_21_n637) );
  INV_X1 p8_mult_21_U648 ( .A(p8_mult_21_n742), .ZN(p8_mult_21_n638) );
  XNOR2_X1 p8_mult_21_U647 ( .A(B2[13]), .B(p8_mult_21_n766), .ZN(
        p8_mult_21_n639) );
  AOI22_X1 p8_mult_21_U646 ( .A1(p8_mult_21_n757), .A2(p8_mult_21_n637), .B1(
        p8_mult_21_n638), .B2(p8_mult_21_n639), .ZN(p8_mult_21_n162) );
  XNOR2_X1 p8_mult_21_U645 ( .A(B2[12]), .B(reg3_reg[11]), .ZN(p8_mult_21_n739) );
  INV_X1 p8_mult_21_U644 ( .A(reg3_reg[9]), .ZN(p8_mult_21_n762) );
  XNOR2_X1 p8_mult_21_U643 ( .A(p8_mult_21_n764), .B(reg3_reg[10]), .ZN(
        p8_mult_21_n774) );
  NAND2_X1 p8_mult_21_U642 ( .A1(p8_mult_21_n725), .A2(p8_mult_21_n774), .ZN(
        p8_mult_21_n727) );
  XNOR2_X1 p8_mult_21_U641 ( .A(B2[13]), .B(reg3_reg[11]), .ZN(p8_mult_21_n741) );
  OAI22_X1 p8_mult_21_U640 ( .A1(p8_mult_21_n739), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n741), .ZN(p8_mult_21_n167) );
  INV_X1 p8_mult_21_U639 ( .A(p8_mult_21_n167), .ZN(p8_mult_21_n168) );
  XNOR2_X1 p8_mult_21_U638 ( .A(B2[12]), .B(reg3_reg[9]), .ZN(p8_mult_21_n722)
         );
  INV_X1 p8_mult_21_U637 ( .A(reg3_reg[7]), .ZN(p8_mult_21_n760) );
  XNOR2_X1 p8_mult_21_U636 ( .A(p8_mult_21_n762), .B(reg3_reg[8]), .ZN(
        p8_mult_21_n773) );
  NAND2_X1 p8_mult_21_U635 ( .A1(p8_mult_21_n708), .A2(p8_mult_21_n773), .ZN(
        p8_mult_21_n710) );
  XNOR2_X1 p8_mult_21_U634 ( .A(B2[13]), .B(reg3_reg[9]), .ZN(p8_mult_21_n724)
         );
  OAI22_X1 p8_mult_21_U633 ( .A1(p8_mult_21_n722), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n724), .ZN(p8_mult_21_n177) );
  INV_X1 p8_mult_21_U632 ( .A(p8_mult_21_n177), .ZN(p8_mult_21_n178) );
  XNOR2_X1 p8_mult_21_U631 ( .A(B2[12]), .B(reg3_reg[7]), .ZN(p8_mult_21_n705)
         );
  INV_X1 p8_mult_21_U630 ( .A(reg3_reg[5]), .ZN(p8_mult_21_n758) );
  XNOR2_X1 p8_mult_21_U629 ( .A(p8_mult_21_n760), .B(reg3_reg[6]), .ZN(
        p8_mult_21_n772) );
  NAND2_X1 p8_mult_21_U628 ( .A1(p8_mult_21_n691), .A2(p8_mult_21_n772), .ZN(
        p8_mult_21_n693) );
  XNOR2_X1 p8_mult_21_U627 ( .A(B2[13]), .B(reg3_reg[7]), .ZN(p8_mult_21_n707)
         );
  OAI22_X1 p8_mult_21_U626 ( .A1(p8_mult_21_n705), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n707), .ZN(p8_mult_21_n191) );
  INV_X1 p8_mult_21_U625 ( .A(p8_mult_21_n191), .ZN(p8_mult_21_n192) );
  XNOR2_X1 p8_mult_21_U624 ( .A(B2[12]), .B(reg3_reg[5]), .ZN(p8_mult_21_n688)
         );
  XNOR2_X1 p8_mult_21_U623 ( .A(p8_mult_21_n758), .B(reg3_reg[4]), .ZN(
        p8_mult_21_n770) );
  NAND2_X1 p8_mult_21_U622 ( .A1(p8_mult_21_n674), .A2(p8_mult_21_n770), .ZN(
        p8_mult_21_n676) );
  XNOR2_X1 p8_mult_21_U621 ( .A(B2[13]), .B(reg3_reg[5]), .ZN(p8_mult_21_n690)
         );
  OAI22_X1 p8_mult_21_U620 ( .A1(p8_mult_21_n688), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n690), .ZN(p8_mult_21_n209) );
  INV_X1 p8_mult_21_U619 ( .A(p8_mult_21_n209), .ZN(p8_mult_21_n210) );
  XNOR2_X1 p8_mult_21_U618 ( .A(B2[12]), .B(reg3_reg[3]), .ZN(p8_mult_21_n670)
         );
  XNOR2_X1 p8_mult_21_U617 ( .A(B2[13]), .B(reg3_reg[3]), .ZN(p8_mult_21_n672)
         );
  OAI22_X1 p8_mult_21_U616 ( .A1(p8_mult_21_n670), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n672), .ZN(p8_mult_21_n231) );
  INV_X1 p8_mult_21_U615 ( .A(p8_mult_21_n231), .ZN(p8_mult_21_n232) );
  XNOR2_X1 p8_mult_21_U614 ( .A(B2[3]), .B(reg3_reg[11]), .ZN(p8_mult_21_n730)
         );
  XNOR2_X1 p8_mult_21_U613 ( .A(B2[4]), .B(reg3_reg[11]), .ZN(p8_mult_21_n731)
         );
  OAI22_X1 p8_mult_21_U612 ( .A1(p8_mult_21_n730), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n731), .ZN(p8_mult_21_n768) );
  XNOR2_X1 p8_mult_21_U611 ( .A(B2[9]), .B(reg3_reg[5]), .ZN(p8_mult_21_n685)
         );
  XNOR2_X1 p8_mult_21_U610 ( .A(B2[10]), .B(reg3_reg[5]), .ZN(p8_mult_21_n686)
         );
  OAI22_X1 p8_mult_21_U609 ( .A1(p8_mult_21_n685), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n686), .ZN(p8_mult_21_n769) );
  OR2_X1 p8_mult_21_U608 ( .A1(p8_mult_21_n768), .A2(p8_mult_21_n769), .ZN(
        p8_mult_21_n243) );
  XNOR2_X1 p8_mult_21_U607 ( .A(p8_mult_21_n768), .B(p8_mult_21_n769), .ZN(
        p8_mult_21_n244) );
  NAND3_X1 p8_mult_21_U606 ( .A1(p8_mult_21_n638), .A2(p8_mult_21_n673), .A3(
        reg3_reg[13]), .ZN(p8_mult_21_n767) );
  OAI21_X1 p8_mult_21_U605 ( .B1(p8_mult_21_n766), .B2(p8_mult_21_n744), .A(
        p8_mult_21_n767), .ZN(p8_mult_21_n317) );
  OR3_X1 p8_mult_21_U604 ( .A1(p8_mult_21_n725), .A2(B2[0]), .A3(
        p8_mult_21_n764), .ZN(p8_mult_21_n765) );
  OAI21_X1 p8_mult_21_U603 ( .B1(p8_mult_21_n764), .B2(p8_mult_21_n727), .A(
        p8_mult_21_n765), .ZN(p8_mult_21_n318) );
  OR3_X1 p8_mult_21_U602 ( .A1(p8_mult_21_n708), .A2(B2[0]), .A3(
        p8_mult_21_n762), .ZN(p8_mult_21_n763) );
  OAI21_X1 p8_mult_21_U601 ( .B1(p8_mult_21_n762), .B2(p8_mult_21_n710), .A(
        p8_mult_21_n763), .ZN(p8_mult_21_n319) );
  OR3_X1 p8_mult_21_U600 ( .A1(p8_mult_21_n691), .A2(B2[0]), .A3(
        p8_mult_21_n760), .ZN(p8_mult_21_n761) );
  OAI21_X1 p8_mult_21_U599 ( .B1(p8_mult_21_n760), .B2(p8_mult_21_n693), .A(
        p8_mult_21_n761), .ZN(p8_mult_21_n320) );
  OR3_X1 p8_mult_21_U598 ( .A1(p8_mult_21_n674), .A2(B2[0]), .A3(
        p8_mult_21_n758), .ZN(p8_mult_21_n759) );
  OAI21_X1 p8_mult_21_U597 ( .B1(p8_mult_21_n758), .B2(p8_mult_21_n676), .A(
        p8_mult_21_n759), .ZN(p8_mult_21_n321) );
  XNOR2_X1 p8_mult_21_U596 ( .A(B2[11]), .B(reg3_reg[13]), .ZN(p8_mult_21_n755) );
  INV_X1 p8_mult_21_U595 ( .A(p8_mult_21_n757), .ZN(p8_mult_21_n756) );
  OAI22_X1 p8_mult_21_U594 ( .A1(p8_mult_21_n755), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n756), .ZN(p8_mult_21_n325) );
  XNOR2_X1 p8_mult_21_U593 ( .A(B2[10]), .B(reg3_reg[13]), .ZN(p8_mult_21_n754) );
  OAI22_X1 p8_mult_21_U592 ( .A1(p8_mult_21_n754), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n755), .ZN(p8_mult_21_n326) );
  XNOR2_X1 p8_mult_21_U591 ( .A(B2[9]), .B(reg3_reg[13]), .ZN(p8_mult_21_n753)
         );
  OAI22_X1 p8_mult_21_U590 ( .A1(p8_mult_21_n753), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n754), .ZN(p8_mult_21_n327) );
  XNOR2_X1 p8_mult_21_U589 ( .A(B2[8]), .B(reg3_reg[13]), .ZN(p8_mult_21_n752)
         );
  OAI22_X1 p8_mult_21_U588 ( .A1(p8_mult_21_n752), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n753), .ZN(p8_mult_21_n328) );
  XNOR2_X1 p8_mult_21_U587 ( .A(B2[7]), .B(reg3_reg[13]), .ZN(p8_mult_21_n751)
         );
  OAI22_X1 p8_mult_21_U586 ( .A1(p8_mult_21_n751), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n752), .ZN(p8_mult_21_n329) );
  XNOR2_X1 p8_mult_21_U585 ( .A(B2[6]), .B(reg3_reg[13]), .ZN(p8_mult_21_n750)
         );
  OAI22_X1 p8_mult_21_U584 ( .A1(p8_mult_21_n750), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n751), .ZN(p8_mult_21_n330) );
  XNOR2_X1 p8_mult_21_U583 ( .A(B2[5]), .B(reg3_reg[13]), .ZN(p8_mult_21_n749)
         );
  OAI22_X1 p8_mult_21_U582 ( .A1(p8_mult_21_n749), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n750), .ZN(p8_mult_21_n331) );
  XNOR2_X1 p8_mult_21_U581 ( .A(B2[4]), .B(reg3_reg[13]), .ZN(p8_mult_21_n748)
         );
  OAI22_X1 p8_mult_21_U580 ( .A1(p8_mult_21_n748), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n749), .ZN(p8_mult_21_n332) );
  XNOR2_X1 p8_mult_21_U579 ( .A(B2[3]), .B(reg3_reg[13]), .ZN(p8_mult_21_n747)
         );
  OAI22_X1 p8_mult_21_U578 ( .A1(p8_mult_21_n747), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n748), .ZN(p8_mult_21_n333) );
  XNOR2_X1 p8_mult_21_U577 ( .A(B2[2]), .B(reg3_reg[13]), .ZN(p8_mult_21_n746)
         );
  OAI22_X1 p8_mult_21_U576 ( .A1(p8_mult_21_n746), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n747), .ZN(p8_mult_21_n334) );
  XNOR2_X1 p8_mult_21_U575 ( .A(B2[1]), .B(reg3_reg[13]), .ZN(p8_mult_21_n745)
         );
  OAI22_X1 p8_mult_21_U574 ( .A1(p8_mult_21_n745), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n746), .ZN(p8_mult_21_n335) );
  XNOR2_X1 p8_mult_21_U573 ( .A(reg3_reg[13]), .B(B2[0]), .ZN(p8_mult_21_n743)
         );
  OAI22_X1 p8_mult_21_U572 ( .A1(p8_mult_21_n743), .A2(p8_mult_21_n744), .B1(
        p8_mult_21_n742), .B2(p8_mult_21_n745), .ZN(p8_mult_21_n336) );
  NOR2_X1 p8_mult_21_U571 ( .A1(p8_mult_21_n673), .A2(p8_mult_21_n742), .ZN(
        p8_mult_21_n337) );
  AOI21_X1 p8_mult_21_U570 ( .B1(p8_mult_21_n727), .B2(p8_mult_21_n725), .A(
        p8_mult_21_n741), .ZN(p8_mult_21_n740) );
  INV_X1 p8_mult_21_U569 ( .A(p8_mult_21_n740), .ZN(p8_mult_21_n338) );
  XNOR2_X1 p8_mult_21_U568 ( .A(B2[11]), .B(reg3_reg[11]), .ZN(p8_mult_21_n738) );
  OAI22_X1 p8_mult_21_U567 ( .A1(p8_mult_21_n738), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n739), .ZN(p8_mult_21_n339) );
  XNOR2_X1 p8_mult_21_U566 ( .A(B2[10]), .B(reg3_reg[11]), .ZN(p8_mult_21_n737) );
  OAI22_X1 p8_mult_21_U565 ( .A1(p8_mult_21_n737), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n738), .ZN(p8_mult_21_n340) );
  XNOR2_X1 p8_mult_21_U564 ( .A(B2[9]), .B(reg3_reg[11]), .ZN(p8_mult_21_n736)
         );
  OAI22_X1 p8_mult_21_U563 ( .A1(p8_mult_21_n736), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n737), .ZN(p8_mult_21_n341) );
  XNOR2_X1 p8_mult_21_U562 ( .A(B2[8]), .B(reg3_reg[11]), .ZN(p8_mult_21_n735)
         );
  OAI22_X1 p8_mult_21_U561 ( .A1(p8_mult_21_n735), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n736), .ZN(p8_mult_21_n342) );
  XNOR2_X1 p8_mult_21_U560 ( .A(B2[7]), .B(reg3_reg[11]), .ZN(p8_mult_21_n734)
         );
  OAI22_X1 p8_mult_21_U559 ( .A1(p8_mult_21_n734), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n735), .ZN(p8_mult_21_n343) );
  XNOR2_X1 p8_mult_21_U558 ( .A(B2[6]), .B(reg3_reg[11]), .ZN(p8_mult_21_n733)
         );
  OAI22_X1 p8_mult_21_U557 ( .A1(p8_mult_21_n733), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n734), .ZN(p8_mult_21_n344) );
  XNOR2_X1 p8_mult_21_U556 ( .A(B2[5]), .B(reg3_reg[11]), .ZN(p8_mult_21_n732)
         );
  OAI22_X1 p8_mult_21_U555 ( .A1(p8_mult_21_n732), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n733), .ZN(p8_mult_21_n345) );
  OAI22_X1 p8_mult_21_U554 ( .A1(p8_mult_21_n731), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n732), .ZN(p8_mult_21_n346) );
  XNOR2_X1 p8_mult_21_U553 ( .A(B2[2]), .B(reg3_reg[11]), .ZN(p8_mult_21_n729)
         );
  OAI22_X1 p8_mult_21_U552 ( .A1(p8_mult_21_n729), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n730), .ZN(p8_mult_21_n348) );
  XNOR2_X1 p8_mult_21_U551 ( .A(B2[1]), .B(reg3_reg[11]), .ZN(p8_mult_21_n728)
         );
  OAI22_X1 p8_mult_21_U550 ( .A1(p8_mult_21_n728), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n729), .ZN(p8_mult_21_n349) );
  XNOR2_X1 p8_mult_21_U549 ( .A(reg3_reg[11]), .B(B2[0]), .ZN(p8_mult_21_n726)
         );
  OAI22_X1 p8_mult_21_U548 ( .A1(p8_mult_21_n726), .A2(p8_mult_21_n727), .B1(
        p8_mult_21_n725), .B2(p8_mult_21_n728), .ZN(p8_mult_21_n350) );
  NOR2_X1 p8_mult_21_U547 ( .A1(p8_mult_21_n673), .A2(p8_mult_21_n725), .ZN(
        p8_mult_21_n351) );
  AOI21_X1 p8_mult_21_U546 ( .B1(p8_mult_21_n710), .B2(p8_mult_21_n708), .A(
        p8_mult_21_n724), .ZN(p8_mult_21_n723) );
  INV_X1 p8_mult_21_U545 ( .A(p8_mult_21_n723), .ZN(p8_mult_21_n352) );
  XNOR2_X1 p8_mult_21_U544 ( .A(B2[11]), .B(reg3_reg[9]), .ZN(p8_mult_21_n721)
         );
  OAI22_X1 p8_mult_21_U543 ( .A1(p8_mult_21_n721), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n722), .ZN(p8_mult_21_n353) );
  XNOR2_X1 p8_mult_21_U542 ( .A(B2[10]), .B(reg3_reg[9]), .ZN(p8_mult_21_n720)
         );
  OAI22_X1 p8_mult_21_U541 ( .A1(p8_mult_21_n720), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n721), .ZN(p8_mult_21_n354) );
  XNOR2_X1 p8_mult_21_U540 ( .A(B2[9]), .B(reg3_reg[9]), .ZN(p8_mult_21_n719)
         );
  OAI22_X1 p8_mult_21_U539 ( .A1(p8_mult_21_n719), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n720), .ZN(p8_mult_21_n355) );
  XNOR2_X1 p8_mult_21_U538 ( .A(B2[8]), .B(reg3_reg[9]), .ZN(p8_mult_21_n718)
         );
  OAI22_X1 p8_mult_21_U537 ( .A1(p8_mult_21_n718), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n719), .ZN(p8_mult_21_n356) );
  XNOR2_X1 p8_mult_21_U536 ( .A(B2[7]), .B(reg3_reg[9]), .ZN(p8_mult_21_n717)
         );
  OAI22_X1 p8_mult_21_U535 ( .A1(p8_mult_21_n717), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n718), .ZN(p8_mult_21_n357) );
  XNOR2_X1 p8_mult_21_U534 ( .A(B2[6]), .B(reg3_reg[9]), .ZN(p8_mult_21_n716)
         );
  OAI22_X1 p8_mult_21_U533 ( .A1(p8_mult_21_n716), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n717), .ZN(p8_mult_21_n358) );
  XNOR2_X1 p8_mult_21_U532 ( .A(B2[5]), .B(reg3_reg[9]), .ZN(p8_mult_21_n715)
         );
  OAI22_X1 p8_mult_21_U531 ( .A1(p8_mult_21_n715), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n716), .ZN(p8_mult_21_n359) );
  XNOR2_X1 p8_mult_21_U530 ( .A(B2[4]), .B(reg3_reg[9]), .ZN(p8_mult_21_n714)
         );
  OAI22_X1 p8_mult_21_U529 ( .A1(p8_mult_21_n714), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n715), .ZN(p8_mult_21_n360) );
  XNOR2_X1 p8_mult_21_U528 ( .A(B2[3]), .B(reg3_reg[9]), .ZN(p8_mult_21_n713)
         );
  OAI22_X1 p8_mult_21_U527 ( .A1(p8_mult_21_n713), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n714), .ZN(p8_mult_21_n361) );
  XNOR2_X1 p8_mult_21_U526 ( .A(B2[2]), .B(reg3_reg[9]), .ZN(p8_mult_21_n712)
         );
  OAI22_X1 p8_mult_21_U525 ( .A1(p8_mult_21_n712), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n713), .ZN(p8_mult_21_n362) );
  XNOR2_X1 p8_mult_21_U524 ( .A(B2[1]), .B(reg3_reg[9]), .ZN(p8_mult_21_n711)
         );
  OAI22_X1 p8_mult_21_U523 ( .A1(p8_mult_21_n711), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n712), .ZN(p8_mult_21_n363) );
  XNOR2_X1 p8_mult_21_U522 ( .A(reg3_reg[9]), .B(B2[0]), .ZN(p8_mult_21_n709)
         );
  OAI22_X1 p8_mult_21_U521 ( .A1(p8_mult_21_n709), .A2(p8_mult_21_n710), .B1(
        p8_mult_21_n708), .B2(p8_mult_21_n711), .ZN(p8_mult_21_n364) );
  NOR2_X1 p8_mult_21_U520 ( .A1(p8_mult_21_n673), .A2(p8_mult_21_n708), .ZN(
        p8_mult_21_n365) );
  AOI21_X1 p8_mult_21_U519 ( .B1(p8_mult_21_n693), .B2(p8_mult_21_n691), .A(
        p8_mult_21_n707), .ZN(p8_mult_21_n706) );
  INV_X1 p8_mult_21_U518 ( .A(p8_mult_21_n706), .ZN(p8_mult_21_n366) );
  XNOR2_X1 p8_mult_21_U517 ( .A(B2[11]), .B(reg3_reg[7]), .ZN(p8_mult_21_n704)
         );
  OAI22_X1 p8_mult_21_U516 ( .A1(p8_mult_21_n704), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n705), .ZN(p8_mult_21_n367) );
  XNOR2_X1 p8_mult_21_U515 ( .A(B2[10]), .B(reg3_reg[7]), .ZN(p8_mult_21_n703)
         );
  OAI22_X1 p8_mult_21_U514 ( .A1(p8_mult_21_n703), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n704), .ZN(p8_mult_21_n368) );
  XNOR2_X1 p8_mult_21_U513 ( .A(B2[9]), .B(reg3_reg[7]), .ZN(p8_mult_21_n702)
         );
  OAI22_X1 p8_mult_21_U512 ( .A1(p8_mult_21_n702), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n703), .ZN(p8_mult_21_n369) );
  XNOR2_X1 p8_mult_21_U511 ( .A(B2[8]), .B(reg3_reg[7]), .ZN(p8_mult_21_n701)
         );
  OAI22_X1 p8_mult_21_U510 ( .A1(p8_mult_21_n701), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n702), .ZN(p8_mult_21_n370) );
  XNOR2_X1 p8_mult_21_U509 ( .A(B2[7]), .B(reg3_reg[7]), .ZN(p8_mult_21_n700)
         );
  OAI22_X1 p8_mult_21_U508 ( .A1(p8_mult_21_n700), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n701), .ZN(p8_mult_21_n371) );
  XNOR2_X1 p8_mult_21_U507 ( .A(B2[6]), .B(reg3_reg[7]), .ZN(p8_mult_21_n699)
         );
  OAI22_X1 p8_mult_21_U506 ( .A1(p8_mult_21_n699), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n700), .ZN(p8_mult_21_n372) );
  XNOR2_X1 p8_mult_21_U505 ( .A(B2[5]), .B(reg3_reg[7]), .ZN(p8_mult_21_n698)
         );
  OAI22_X1 p8_mult_21_U504 ( .A1(p8_mult_21_n698), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n699), .ZN(p8_mult_21_n373) );
  XNOR2_X1 p8_mult_21_U503 ( .A(B2[4]), .B(reg3_reg[7]), .ZN(p8_mult_21_n697)
         );
  OAI22_X1 p8_mult_21_U502 ( .A1(p8_mult_21_n697), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n698), .ZN(p8_mult_21_n374) );
  XNOR2_X1 p8_mult_21_U501 ( .A(B2[3]), .B(reg3_reg[7]), .ZN(p8_mult_21_n696)
         );
  OAI22_X1 p8_mult_21_U500 ( .A1(p8_mult_21_n696), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n697), .ZN(p8_mult_21_n375) );
  XNOR2_X1 p8_mult_21_U499 ( .A(B2[2]), .B(reg3_reg[7]), .ZN(p8_mult_21_n695)
         );
  OAI22_X1 p8_mult_21_U498 ( .A1(p8_mult_21_n695), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n696), .ZN(p8_mult_21_n376) );
  XNOR2_X1 p8_mult_21_U497 ( .A(B2[1]), .B(reg3_reg[7]), .ZN(p8_mult_21_n694)
         );
  OAI22_X1 p8_mult_21_U496 ( .A1(p8_mult_21_n694), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n695), .ZN(p8_mult_21_n377) );
  XNOR2_X1 p8_mult_21_U495 ( .A(reg3_reg[7]), .B(B2[0]), .ZN(p8_mult_21_n692)
         );
  OAI22_X1 p8_mult_21_U494 ( .A1(p8_mult_21_n692), .A2(p8_mult_21_n693), .B1(
        p8_mult_21_n691), .B2(p8_mult_21_n694), .ZN(p8_mult_21_n378) );
  NOR2_X1 p8_mult_21_U493 ( .A1(p8_mult_21_n673), .A2(p8_mult_21_n691), .ZN(
        p8_mult_21_n379) );
  AOI21_X1 p8_mult_21_U492 ( .B1(p8_mult_21_n676), .B2(p8_mult_21_n674), .A(
        p8_mult_21_n690), .ZN(p8_mult_21_n689) );
  INV_X1 p8_mult_21_U491 ( .A(p8_mult_21_n689), .ZN(p8_mult_21_n380) );
  XNOR2_X1 p8_mult_21_U490 ( .A(B2[11]), .B(reg3_reg[5]), .ZN(p8_mult_21_n687)
         );
  OAI22_X1 p8_mult_21_U489 ( .A1(p8_mult_21_n687), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n688), .ZN(p8_mult_21_n381) );
  OAI22_X1 p8_mult_21_U488 ( .A1(p8_mult_21_n686), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n687), .ZN(p8_mult_21_n382) );
  XNOR2_X1 p8_mult_21_U487 ( .A(B2[8]), .B(reg3_reg[5]), .ZN(p8_mult_21_n684)
         );
  OAI22_X1 p8_mult_21_U486 ( .A1(p8_mult_21_n684), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n685), .ZN(p8_mult_21_n384) );
  XNOR2_X1 p8_mult_21_U485 ( .A(B2[7]), .B(reg3_reg[5]), .ZN(p8_mult_21_n683)
         );
  OAI22_X1 p8_mult_21_U484 ( .A1(p8_mult_21_n683), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n684), .ZN(p8_mult_21_n385) );
  XNOR2_X1 p8_mult_21_U483 ( .A(B2[6]), .B(reg3_reg[5]), .ZN(p8_mult_21_n682)
         );
  OAI22_X1 p8_mult_21_U482 ( .A1(p8_mult_21_n682), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n683), .ZN(p8_mult_21_n386) );
  XNOR2_X1 p8_mult_21_U481 ( .A(B2[5]), .B(reg3_reg[5]), .ZN(p8_mult_21_n681)
         );
  OAI22_X1 p8_mult_21_U480 ( .A1(p8_mult_21_n681), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n682), .ZN(p8_mult_21_n387) );
  XNOR2_X1 p8_mult_21_U479 ( .A(B2[4]), .B(reg3_reg[5]), .ZN(p8_mult_21_n680)
         );
  OAI22_X1 p8_mult_21_U478 ( .A1(p8_mult_21_n680), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n681), .ZN(p8_mult_21_n388) );
  XNOR2_X1 p8_mult_21_U477 ( .A(B2[3]), .B(reg3_reg[5]), .ZN(p8_mult_21_n679)
         );
  OAI22_X1 p8_mult_21_U476 ( .A1(p8_mult_21_n679), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n680), .ZN(p8_mult_21_n389) );
  XNOR2_X1 p8_mult_21_U475 ( .A(B2[2]), .B(reg3_reg[5]), .ZN(p8_mult_21_n678)
         );
  OAI22_X1 p8_mult_21_U474 ( .A1(p8_mult_21_n678), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n679), .ZN(p8_mult_21_n390) );
  XNOR2_X1 p8_mult_21_U473 ( .A(B2[1]), .B(reg3_reg[5]), .ZN(p8_mult_21_n677)
         );
  OAI22_X1 p8_mult_21_U472 ( .A1(p8_mult_21_n677), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n678), .ZN(p8_mult_21_n391) );
  XNOR2_X1 p8_mult_21_U471 ( .A(reg3_reg[5]), .B(B2[0]), .ZN(p8_mult_21_n675)
         );
  OAI22_X1 p8_mult_21_U470 ( .A1(p8_mult_21_n675), .A2(p8_mult_21_n676), .B1(
        p8_mult_21_n674), .B2(p8_mult_21_n677), .ZN(p8_mult_21_n392) );
  NOR2_X1 p8_mult_21_U469 ( .A1(p8_mult_21_n673), .A2(p8_mult_21_n674), .ZN(
        p8_mult_21_n393) );
  AOI21_X1 p8_mult_21_U468 ( .B1(p8_mult_21_n657), .B2(p8_mult_21_n658), .A(
        p8_mult_21_n672), .ZN(p8_mult_21_n671) );
  INV_X1 p8_mult_21_U467 ( .A(p8_mult_21_n671), .ZN(p8_mult_21_n394) );
  XNOR2_X1 p8_mult_21_U466 ( .A(B2[11]), .B(reg3_reg[3]), .ZN(p8_mult_21_n669)
         );
  OAI22_X1 p8_mult_21_U465 ( .A1(p8_mult_21_n669), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n670), .ZN(p8_mult_21_n395) );
  XNOR2_X1 p8_mult_21_U464 ( .A(B2[10]), .B(reg3_reg[3]), .ZN(p8_mult_21_n668)
         );
  OAI22_X1 p8_mult_21_U463 ( .A1(p8_mult_21_n668), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n669), .ZN(p8_mult_21_n396) );
  XNOR2_X1 p8_mult_21_U462 ( .A(B2[9]), .B(reg3_reg[3]), .ZN(p8_mult_21_n667)
         );
  OAI22_X1 p8_mult_21_U461 ( .A1(p8_mult_21_n667), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n668), .ZN(p8_mult_21_n397) );
  XNOR2_X1 p8_mult_21_U460 ( .A(B2[8]), .B(reg3_reg[3]), .ZN(p8_mult_21_n666)
         );
  OAI22_X1 p8_mult_21_U459 ( .A1(p8_mult_21_n666), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n667), .ZN(p8_mult_21_n398) );
  XNOR2_X1 p8_mult_21_U458 ( .A(B2[7]), .B(reg3_reg[3]), .ZN(p8_mult_21_n665)
         );
  OAI22_X1 p8_mult_21_U457 ( .A1(p8_mult_21_n665), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n666), .ZN(p8_mult_21_n399) );
  XNOR2_X1 p8_mult_21_U456 ( .A(B2[6]), .B(reg3_reg[3]), .ZN(p8_mult_21_n664)
         );
  OAI22_X1 p8_mult_21_U455 ( .A1(p8_mult_21_n664), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n665), .ZN(p8_mult_21_n400) );
  XNOR2_X1 p8_mult_21_U454 ( .A(B2[5]), .B(reg3_reg[3]), .ZN(p8_mult_21_n663)
         );
  OAI22_X1 p8_mult_21_U453 ( .A1(p8_mult_21_n663), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n664), .ZN(p8_mult_21_n401) );
  XNOR2_X1 p8_mult_21_U452 ( .A(B2[4]), .B(reg3_reg[3]), .ZN(p8_mult_21_n662)
         );
  OAI22_X1 p8_mult_21_U451 ( .A1(p8_mult_21_n662), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n663), .ZN(p8_mult_21_n402) );
  XNOR2_X1 p8_mult_21_U450 ( .A(B2[3]), .B(reg3_reg[3]), .ZN(p8_mult_21_n661)
         );
  OAI22_X1 p8_mult_21_U449 ( .A1(p8_mult_21_n661), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n662), .ZN(p8_mult_21_n403) );
  XNOR2_X1 p8_mult_21_U448 ( .A(B2[2]), .B(reg3_reg[3]), .ZN(p8_mult_21_n660)
         );
  OAI22_X1 p8_mult_21_U447 ( .A1(p8_mult_21_n660), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n661), .ZN(p8_mult_21_n404) );
  XNOR2_X1 p8_mult_21_U446 ( .A(B2[1]), .B(reg3_reg[3]), .ZN(p8_mult_21_n659)
         );
  OAI22_X1 p8_mult_21_U445 ( .A1(p8_mult_21_n659), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n660), .ZN(p8_mult_21_n405) );
  XNOR2_X1 p8_mult_21_U444 ( .A(reg3_reg[3]), .B(B2[0]), .ZN(p8_mult_21_n656)
         );
  OAI22_X1 p8_mult_21_U443 ( .A1(p8_mult_21_n656), .A2(p8_mult_21_n657), .B1(
        p8_mult_21_n658), .B2(p8_mult_21_n659), .ZN(p8_mult_21_n406) );
  XOR2_X1 p8_mult_21_U442 ( .A(B2[13]), .B(p8_mult_21_n655), .Z(
        p8_mult_21_n653) );
  AOI21_X1 p8_mult_21_U441 ( .B1(p8_mult_21_n641), .B2(p8_mult_21_n643), .A(
        p8_mult_21_n653), .ZN(p8_mult_21_n654) );
  INV_X1 p8_mult_21_U440 ( .A(p8_mult_21_n654), .ZN(p8_mult_21_n408) );
  XNOR2_X1 p8_mult_21_U439 ( .A(B2[12]), .B(reg3_reg[1]), .ZN(p8_mult_21_n652)
         );
  OAI22_X1 p8_mult_21_U438 ( .A1(p8_mult_21_n652), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n653), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n409) );
  XNOR2_X1 p8_mult_21_U437 ( .A(B2[11]), .B(reg3_reg[1]), .ZN(p8_mult_21_n651)
         );
  OAI22_X1 p8_mult_21_U436 ( .A1(p8_mult_21_n651), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n652), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n410) );
  XNOR2_X1 p8_mult_21_U435 ( .A(B2[10]), .B(reg3_reg[1]), .ZN(p8_mult_21_n650)
         );
  OAI22_X1 p8_mult_21_U434 ( .A1(p8_mult_21_n650), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n651), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n411) );
  XNOR2_X1 p8_mult_21_U433 ( .A(B2[9]), .B(reg3_reg[1]), .ZN(p8_mult_21_n649)
         );
  OAI22_X1 p8_mult_21_U432 ( .A1(p8_mult_21_n649), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n650), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n412) );
  XNOR2_X1 p8_mult_21_U431 ( .A(B2[8]), .B(reg3_reg[1]), .ZN(p8_mult_21_n648)
         );
  OAI22_X1 p8_mult_21_U430 ( .A1(p8_mult_21_n648), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n649), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n413) );
  XNOR2_X1 p8_mult_21_U429 ( .A(B2[7]), .B(reg3_reg[1]), .ZN(p8_mult_21_n647)
         );
  OAI22_X1 p8_mult_21_U428 ( .A1(p8_mult_21_n647), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n648), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n414) );
  XNOR2_X1 p8_mult_21_U427 ( .A(B2[6]), .B(reg3_reg[1]), .ZN(p8_mult_21_n646)
         );
  OAI22_X1 p8_mult_21_U426 ( .A1(p8_mult_21_n646), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n647), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n415) );
  XNOR2_X1 p8_mult_21_U425 ( .A(B2[5]), .B(reg3_reg[1]), .ZN(p8_mult_21_n645)
         );
  OAI22_X1 p8_mult_21_U424 ( .A1(p8_mult_21_n645), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n646), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n416) );
  XNOR2_X1 p8_mult_21_U423 ( .A(B2[4]), .B(reg3_reg[1]), .ZN(p8_mult_21_n644)
         );
  OAI22_X1 p8_mult_21_U422 ( .A1(p8_mult_21_n644), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n645), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n417) );
  XNOR2_X1 p8_mult_21_U421 ( .A(B2[3]), .B(reg3_reg[1]), .ZN(p8_mult_21_n642)
         );
  OAI22_X1 p8_mult_21_U420 ( .A1(p8_mult_21_n642), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n644), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n418) );
  OAI22_X1 p8_mult_21_U419 ( .A1(p8_mult_21_n640), .A2(p8_mult_21_n641), .B1(
        p8_mult_21_n642), .B2(p8_mult_21_n643), .ZN(p8_mult_21_n419) );
  OAI21_X1 p8_mult_21_U418 ( .B1(p8_mult_21_n637), .B2(p8_mult_21_n638), .A(
        p8_mult_21_n639), .ZN(p8_mult_21_n636) );
  XOR2_X1 p8_mult_21_U417 ( .A(p8_mult_21_n636), .B(p8_mult_21_n136), .Z(
        p8_mult_21_n635) );
  XNOR2_X1 p8_mult_21_U416 ( .A(p8_mult_21_n162), .B(p8_mult_21_n635), .ZN(
        temp3[13]) );
  XOR2_X2 p8_mult_21_U415 ( .A(reg3_reg[12]), .B(p8_mult_21_n764), .Z(
        p8_mult_21_n742) );
  XOR2_X2 p8_mult_21_U414 ( .A(reg3_reg[10]), .B(p8_mult_21_n762), .Z(
        p8_mult_21_n725) );
  XOR2_X2 p8_mult_21_U413 ( .A(reg3_reg[8]), .B(p8_mult_21_n760), .Z(
        p8_mult_21_n708) );
  XOR2_X2 p8_mult_21_U412 ( .A(reg3_reg[6]), .B(p8_mult_21_n758), .Z(
        p8_mult_21_n691) );
  XOR2_X2 p8_mult_21_U411 ( .A(reg3_reg[4]), .B(p8_mult_21_n771), .Z(
        p8_mult_21_n674) );
  INV_X1 p8_mult_21_U410 ( .A(reg3_reg[0]), .ZN(p8_mult_21_n643) );
  INV_X1 p8_mult_21_U409 ( .A(p8_mult_21_n798), .ZN(p8_mult_21_n658) );
  HA_X1 p8_mult_21_U145 ( .A(p8_mult_21_n406), .B(p8_mult_21_n419), .CO(
        p8_mult_21_n315), .S(p8_mult_21_n316) );
  FA_X1 p8_mult_21_U144 ( .A(p8_mult_21_n418), .B(p8_mult_21_n393), .CI(
        p8_mult_21_n405), .CO(p8_mult_21_n313), .S(p8_mult_21_n314) );
  HA_X1 p8_mult_21_U143 ( .A(p8_mult_21_n321), .B(p8_mult_21_n392), .CO(
        p8_mult_21_n311), .S(p8_mult_21_n312) );
  FA_X1 p8_mult_21_U142 ( .A(p8_mult_21_n404), .B(p8_mult_21_n417), .CI(
        p8_mult_21_n312), .CO(p8_mult_21_n309), .S(p8_mult_21_n310) );
  FA_X1 p8_mult_21_U141 ( .A(p8_mult_21_n416), .B(p8_mult_21_n379), .CI(
        p8_mult_21_n403), .CO(p8_mult_21_n307), .S(p8_mult_21_n308) );
  FA_X1 p8_mult_21_U140 ( .A(p8_mult_21_n311), .B(p8_mult_21_n391), .CI(
        p8_mult_21_n308), .CO(p8_mult_21_n305), .S(p8_mult_21_n306) );
  HA_X1 p8_mult_21_U139 ( .A(p8_mult_21_n320), .B(p8_mult_21_n378), .CO(
        p8_mult_21_n303), .S(p8_mult_21_n304) );
  FA_X1 p8_mult_21_U138 ( .A(p8_mult_21_n390), .B(p8_mult_21_n415), .CI(
        p8_mult_21_n402), .CO(p8_mult_21_n301), .S(p8_mult_21_n302) );
  FA_X1 p8_mult_21_U137 ( .A(p8_mult_21_n307), .B(p8_mult_21_n304), .CI(
        p8_mult_21_n302), .CO(p8_mult_21_n299), .S(p8_mult_21_n300) );
  FA_X1 p8_mult_21_U136 ( .A(p8_mult_21_n389), .B(p8_mult_21_n365), .CI(
        p8_mult_21_n414), .CO(p8_mult_21_n297), .S(p8_mult_21_n298) );
  FA_X1 p8_mult_21_U135 ( .A(p8_mult_21_n377), .B(p8_mult_21_n401), .CI(
        p8_mult_21_n303), .CO(p8_mult_21_n295), .S(p8_mult_21_n296) );
  FA_X1 p8_mult_21_U134 ( .A(p8_mult_21_n298), .B(p8_mult_21_n301), .CI(
        p8_mult_21_n296), .CO(p8_mult_21_n293), .S(p8_mult_21_n294) );
  HA_X1 p8_mult_21_U133 ( .A(p8_mult_21_n319), .B(p8_mult_21_n364), .CO(
        p8_mult_21_n291), .S(p8_mult_21_n292) );
  FA_X1 p8_mult_21_U132 ( .A(p8_mult_21_n376), .B(p8_mult_21_n388), .CI(
        p8_mult_21_n400), .CO(p8_mult_21_n289), .S(p8_mult_21_n290) );
  FA_X1 p8_mult_21_U131 ( .A(p8_mult_21_n292), .B(p8_mult_21_n413), .CI(
        p8_mult_21_n297), .CO(p8_mult_21_n287), .S(p8_mult_21_n288) );
  FA_X1 p8_mult_21_U130 ( .A(p8_mult_21_n290), .B(p8_mult_21_n295), .CI(
        p8_mult_21_n288), .CO(p8_mult_21_n285), .S(p8_mult_21_n286) );
  FA_X1 p8_mult_21_U129 ( .A(p8_mult_21_n375), .B(p8_mult_21_n351), .CI(
        p8_mult_21_n412), .CO(p8_mult_21_n283), .S(p8_mult_21_n284) );
  FA_X1 p8_mult_21_U128 ( .A(p8_mult_21_n363), .B(p8_mult_21_n399), .CI(
        p8_mult_21_n387), .CO(p8_mult_21_n281), .S(p8_mult_21_n282) );
  FA_X1 p8_mult_21_U127 ( .A(p8_mult_21_n289), .B(p8_mult_21_n291), .CI(
        p8_mult_21_n284), .CO(p8_mult_21_n279), .S(p8_mult_21_n280) );
  FA_X1 p8_mult_21_U126 ( .A(p8_mult_21_n287), .B(p8_mult_21_n282), .CI(
        p8_mult_21_n280), .CO(p8_mult_21_n277), .S(p8_mult_21_n278) );
  HA_X1 p8_mult_21_U125 ( .A(p8_mult_21_n318), .B(p8_mult_21_n350), .CO(
        p8_mult_21_n275), .S(p8_mult_21_n276) );
  FA_X1 p8_mult_21_U124 ( .A(p8_mult_21_n362), .B(p8_mult_21_n386), .CI(
        p8_mult_21_n411), .CO(p8_mult_21_n273), .S(p8_mult_21_n274) );
  FA_X1 p8_mult_21_U123 ( .A(p8_mult_21_n374), .B(p8_mult_21_n398), .CI(
        p8_mult_21_n276), .CO(p8_mult_21_n271), .S(p8_mult_21_n272) );
  FA_X1 p8_mult_21_U122 ( .A(p8_mult_21_n281), .B(p8_mult_21_n283), .CI(
        p8_mult_21_n274), .CO(p8_mult_21_n269), .S(p8_mult_21_n270) );
  FA_X1 p8_mult_21_U121 ( .A(p8_mult_21_n279), .B(p8_mult_21_n272), .CI(
        p8_mult_21_n270), .CO(p8_mult_21_n267), .S(p8_mult_21_n268) );
  FA_X1 p8_mult_21_U120 ( .A(p8_mult_21_n361), .B(p8_mult_21_n337), .CI(
        p8_mult_21_n410), .CO(p8_mult_21_n265), .S(p8_mult_21_n266) );
  FA_X1 p8_mult_21_U109 ( .A(p8_mult_21_n349), .B(p8_mult_21_n397), .CI(
        p8_mult_21_n373), .CO(p8_mult_21_n263), .S(p8_mult_21_n264) );
  FA_X1 p8_mult_21_U108 ( .A(p8_mult_21_n275), .B(p8_mult_21_n385), .CI(
        p8_mult_21_n273), .CO(p8_mult_21_n261), .S(p8_mult_21_n262) );
  FA_X1 p8_mult_21_U107 ( .A(p8_mult_21_n264), .B(p8_mult_21_n266), .CI(
        p8_mult_21_n271), .CO(p8_mult_21_n259), .S(p8_mult_21_n260) );
  FA_X1 p8_mult_21_U106 ( .A(p8_mult_21_n262), .B(p8_mult_21_n269), .CI(
        p8_mult_21_n260), .CO(p8_mult_21_n257), .S(p8_mult_21_n258) );
  HA_X1 p8_mult_21_U105 ( .A(p8_mult_21_n317), .B(p8_mult_21_n336), .CO(
        p8_mult_21_n255), .S(p8_mult_21_n256) );
  FA_X1 p8_mult_21_U104 ( .A(p8_mult_21_n409), .B(p8_mult_21_n372), .CI(
        p8_mult_21_n396), .CO(p8_mult_21_n253), .S(p8_mult_21_n254) );
  FA_X1 p8_mult_21_U103 ( .A(p8_mult_21_n348), .B(p8_mult_21_n384), .CI(
        p8_mult_21_n360), .CO(p8_mult_21_n251), .S(p8_mult_21_n252) );
  FA_X1 p8_mult_21_U102 ( .A(p8_mult_21_n265), .B(p8_mult_21_n256), .CI(
        p8_mult_21_n263), .CO(p8_mult_21_n249), .S(p8_mult_21_n250) );
  FA_X1 p8_mult_21_U101 ( .A(p8_mult_21_n254), .B(p8_mult_21_n252), .CI(
        p8_mult_21_n261), .CO(p8_mult_21_n247), .S(p8_mult_21_n248) );
  FA_X1 p8_mult_21_U100 ( .A(p8_mult_21_n259), .B(p8_mult_21_n250), .CI(
        p8_mult_21_n248), .CO(p8_mult_21_n245), .S(p8_mult_21_n246) );
  FA_X1 p8_mult_21_U97 ( .A(p8_mult_21_n395), .B(p8_mult_21_n359), .CI(
        p8_mult_21_n408), .CO(p8_mult_21_n241), .S(p8_mult_21_n242) );
  FA_X1 p8_mult_21_U96 ( .A(p8_mult_21_n335), .B(p8_mult_21_n371), .CI(
        p8_mult_21_n255), .CO(p8_mult_21_n239), .S(p8_mult_21_n240) );
  FA_X1 p8_mult_21_U95 ( .A(p8_mult_21_n253), .B(p8_mult_21_n244), .CI(
        p8_mult_21_n251), .CO(p8_mult_21_n237), .S(p8_mult_21_n238) );
  FA_X1 p8_mult_21_U94 ( .A(p8_mult_21_n240), .B(p8_mult_21_n242), .CI(
        p8_mult_21_n249), .CO(p8_mult_21_n235), .S(p8_mult_21_n236) );
  FA_X1 p8_mult_21_U93 ( .A(p8_mult_21_n247), .B(p8_mult_21_n238), .CI(
        p8_mult_21_n236), .CO(p8_mult_21_n233), .S(p8_mult_21_n234) );
  FA_X1 p8_mult_21_U91 ( .A(p8_mult_21_n382), .B(p8_mult_21_n346), .CI(
        p8_mult_21_n232), .CO(p8_mult_21_n229), .S(p8_mult_21_n230) );
  FA_X1 p8_mult_21_U90 ( .A(p8_mult_21_n334), .B(p8_mult_21_n370), .CI(
        p8_mult_21_n358), .CO(p8_mult_21_n227), .S(p8_mult_21_n228) );
  FA_X1 p8_mult_21_U89 ( .A(p8_mult_21_n241), .B(p8_mult_21_n243), .CI(
        p8_mult_21_n239), .CO(p8_mult_21_n225), .S(p8_mult_21_n226) );
  FA_X1 p8_mult_21_U88 ( .A(p8_mult_21_n230), .B(p8_mult_21_n228), .CI(
        p8_mult_21_n237), .CO(p8_mult_21_n223), .S(p8_mult_21_n224) );
  FA_X1 p8_mult_21_U87 ( .A(p8_mult_21_n235), .B(p8_mult_21_n226), .CI(
        p8_mult_21_n224), .CO(p8_mult_21_n221), .S(p8_mult_21_n222) );
  FA_X1 p8_mult_21_U86 ( .A(p8_mult_21_n231), .B(p8_mult_21_n333), .CI(
        p8_mult_21_n394), .CO(p8_mult_21_n219), .S(p8_mult_21_n220) );
  FA_X1 p8_mult_21_U85 ( .A(p8_mult_21_n345), .B(p8_mult_21_n381), .CI(
        p8_mult_21_n357), .CO(p8_mult_21_n217), .S(p8_mult_21_n218) );
  FA_X1 p8_mult_21_U84 ( .A(p8_mult_21_n229), .B(p8_mult_21_n369), .CI(
        p8_mult_21_n227), .CO(p8_mult_21_n215), .S(p8_mult_21_n216) );
  FA_X1 p8_mult_21_U83 ( .A(p8_mult_21_n220), .B(p8_mult_21_n218), .CI(
        p8_mult_21_n225), .CO(p8_mult_21_n213), .S(p8_mult_21_n214) );
  FA_X1 p8_mult_21_U82 ( .A(p8_mult_21_n223), .B(p8_mult_21_n216), .CI(
        p8_mult_21_n214), .CO(p8_mult_21_n211), .S(p8_mult_21_n212) );
  FA_X1 p8_mult_21_U80 ( .A(p8_mult_21_n368), .B(p8_mult_21_n344), .CI(
        p8_mult_21_n210), .CO(p8_mult_21_n207), .S(p8_mult_21_n208) );
  FA_X1 p8_mult_21_U79 ( .A(p8_mult_21_n332), .B(p8_mult_21_n356), .CI(
        p8_mult_21_n219), .CO(p8_mult_21_n205), .S(p8_mult_21_n206) );
  FA_X1 p8_mult_21_U78 ( .A(p8_mult_21_n208), .B(p8_mult_21_n217), .CI(
        p8_mult_21_n215), .CO(p8_mult_21_n203), .S(p8_mult_21_n204) );
  FA_X1 p8_mult_21_U77 ( .A(p8_mult_21_n213), .B(p8_mult_21_n206), .CI(
        p8_mult_21_n204), .CO(p8_mult_21_n201), .S(p8_mult_21_n202) );
  FA_X1 p8_mult_21_U76 ( .A(p8_mult_21_n209), .B(p8_mult_21_n331), .CI(
        p8_mult_21_n380), .CO(p8_mult_21_n199), .S(p8_mult_21_n200) );
  FA_X1 p8_mult_21_U75 ( .A(p8_mult_21_n355), .B(p8_mult_21_n343), .CI(
        p8_mult_21_n367), .CO(p8_mult_21_n197), .S(p8_mult_21_n198) );
  FA_X1 p8_mult_21_U74 ( .A(p8_mult_21_n198), .B(p8_mult_21_n207), .CI(
        p8_mult_21_n200), .CO(p8_mult_21_n195), .S(p8_mult_21_n196) );
  FA_X1 p8_mult_21_U73 ( .A(p8_mult_21_n203), .B(p8_mult_21_n205), .CI(
        p8_mult_21_n196), .CO(p8_mult_21_n193), .S(p8_mult_21_n194) );
  FA_X1 p8_mult_21_U71 ( .A(p8_mult_21_n330), .B(p8_mult_21_n342), .CI(
        p8_mult_21_n192), .CO(p8_mult_21_n189), .S(p8_mult_21_n190) );
  FA_X1 p8_mult_21_U70 ( .A(p8_mult_21_n199), .B(p8_mult_21_n354), .CI(
        p8_mult_21_n197), .CO(p8_mult_21_n187), .S(p8_mult_21_n188) );
  FA_X1 p8_mult_21_U69 ( .A(p8_mult_21_n188), .B(p8_mult_21_n190), .CI(
        p8_mult_21_n195), .CO(p8_mult_21_n185), .S(p8_mult_21_n186) );
  FA_X1 p8_mult_21_U68 ( .A(p8_mult_21_n191), .B(p8_mult_21_n329), .CI(
        p8_mult_21_n366), .CO(p8_mult_21_n183), .S(p8_mult_21_n184) );
  FA_X1 p8_mult_21_U67 ( .A(p8_mult_21_n341), .B(p8_mult_21_n353), .CI(
        p8_mult_21_n189), .CO(p8_mult_21_n181), .S(p8_mult_21_n182) );
  FA_X1 p8_mult_21_U66 ( .A(p8_mult_21_n187), .B(p8_mult_21_n184), .CI(
        p8_mult_21_n182), .CO(p8_mult_21_n179), .S(p8_mult_21_n180) );
  FA_X1 p8_mult_21_U64 ( .A(p8_mult_21_n328), .B(p8_mult_21_n340), .CI(
        p8_mult_21_n178), .CO(p8_mult_21_n175), .S(p8_mult_21_n176) );
  FA_X1 p8_mult_21_U63 ( .A(p8_mult_21_n176), .B(p8_mult_21_n183), .CI(
        p8_mult_21_n181), .CO(p8_mult_21_n173), .S(p8_mult_21_n174) );
  FA_X1 p8_mult_21_U62 ( .A(p8_mult_21_n327), .B(p8_mult_21_n177), .CI(
        p8_mult_21_n352), .CO(p8_mult_21_n171), .S(p8_mult_21_n172) );
  FA_X1 p8_mult_21_U61 ( .A(p8_mult_21_n175), .B(p8_mult_21_n339), .CI(
        p8_mult_21_n172), .CO(p8_mult_21_n169), .S(p8_mult_21_n170) );
  FA_X1 p8_mult_21_U59 ( .A(p8_mult_21_n168), .B(p8_mult_21_n326), .CI(
        p8_mult_21_n171), .CO(p8_mult_21_n165), .S(p8_mult_21_n166) );
  FA_X1 p8_mult_21_U58 ( .A(p8_mult_21_n325), .B(p8_mult_21_n167), .CI(
        p8_mult_21_n338), .CO(p8_mult_21_n163), .S(p8_mult_21_n164) );
  FA_X1 p8_mult_21_U44 ( .A(p8_mult_21_n246), .B(p8_mult_21_n257), .CI(
        p8_mult_21_n149), .CO(p8_mult_21_n148), .S(temp3[0]) );
  FA_X1 p8_mult_21_U43 ( .A(p8_mult_21_n234), .B(p8_mult_21_n245), .CI(
        p8_mult_21_n148), .CO(p8_mult_21_n147), .S(temp3[1]) );
  FA_X1 p8_mult_21_U42 ( .A(p8_mult_21_n222), .B(p8_mult_21_n233), .CI(
        p8_mult_21_n147), .CO(p8_mult_21_n146), .S(temp3[2]) );
  FA_X1 p8_mult_21_U41 ( .A(p8_mult_21_n212), .B(p8_mult_21_n221), .CI(
        p8_mult_21_n146), .CO(p8_mult_21_n145), .S(temp3[3]) );
  FA_X1 p8_mult_21_U40 ( .A(p8_mult_21_n202), .B(p8_mult_21_n211), .CI(
        p8_mult_21_n145), .CO(p8_mult_21_n144), .S(temp3[4]) );
  FA_X1 p8_mult_21_U39 ( .A(p8_mult_21_n194), .B(p8_mult_21_n201), .CI(
        p8_mult_21_n144), .CO(p8_mult_21_n143), .S(temp3[5]) );
  FA_X1 p8_mult_21_U38 ( .A(p8_mult_21_n186), .B(p8_mult_21_n193), .CI(
        p8_mult_21_n143), .CO(p8_mult_21_n142), .S(temp3[6]) );
  FA_X1 p8_mult_21_U37 ( .A(p8_mult_21_n180), .B(p8_mult_21_n185), .CI(
        p8_mult_21_n142), .CO(p8_mult_21_n141), .S(temp3[7]) );
  FA_X1 p8_mult_21_U30 ( .A(p8_mult_21_n174), .B(p8_mult_21_n179), .CI(
        p8_mult_21_n141), .CO(p8_mult_21_n140), .S(temp3[8]) );
  FA_X1 p8_mult_21_U20 ( .A(p8_mult_21_n170), .B(p8_mult_21_n173), .CI(
        p8_mult_21_n140), .CO(p8_mult_21_n139), .S(temp3[9]) );
  FA_X1 p8_mult_21_U10 ( .A(p8_mult_21_n166), .B(p8_mult_21_n169), .CI(
        p8_mult_21_n139), .CO(p8_mult_21_n138), .S(temp3[10]) );
  FA_X1 p8_mult_21_U9 ( .A(p8_mult_21_n165), .B(p8_mult_21_n164), .CI(
        p8_mult_21_n138), .CO(p8_mult_21_n137), .S(temp3[11]) );
  FA_X1 p8_mult_21_U8 ( .A(p8_mult_21_n163), .B(p8_mult_21_n162), .CI(
        p8_mult_21_n137), .CO(p8_mult_21_n136), .S(temp3[12]) );
  NAND2_X1 REG3_1_U34 ( .A1(temp3[4]), .A2(REG3_1_n43), .ZN(REG3_1_n85) );
  OAI21_X1 REG3_1_U33 ( .B1(REG3_1_n45), .B2(REG3_1_n66), .A(REG3_1_n85), .ZN(
        REG3_1_n57) );
  NAND2_X1 REG3_1_U32 ( .A1(temp3[3]), .A2(REG3_1_n43), .ZN(REG3_1_n86) );
  OAI21_X1 REG3_1_U31 ( .B1(REG3_1_n45), .B2(REG3_1_n65), .A(REG3_1_n86), .ZN(
        REG3_1_n58) );
  NAND2_X1 REG3_1_U30 ( .A1(temp3[2]), .A2(REG3_1_n43), .ZN(REG3_1_n87) );
  OAI21_X1 REG3_1_U29 ( .B1(REG3_1_n45), .B2(REG3_1_n64), .A(REG3_1_n87), .ZN(
        REG3_1_n59) );
  NAND2_X1 REG3_1_U28 ( .A1(temp3[5]), .A2(REG3_1_n43), .ZN(REG3_1_n84) );
  OAI21_X1 REG3_1_U27 ( .B1(REG3_1_n44), .B2(REG3_1_n67), .A(REG3_1_n84), .ZN(
        REG3_1_n56) );
  NAND2_X1 REG3_1_U26 ( .A1(temp3[9]), .A2(REG3_1_n43), .ZN(REG3_1_n80) );
  OAI21_X1 REG3_1_U25 ( .B1(REG3_1_n44), .B2(REG3_1_n71), .A(REG3_1_n80), .ZN(
        REG3_1_n52) );
  NAND2_X1 REG3_1_U24 ( .A1(temp3[8]), .A2(REG3_1_n44), .ZN(REG3_1_n81) );
  OAI21_X1 REG3_1_U23 ( .B1(REG3_1_n44), .B2(REG3_1_n70), .A(REG3_1_n81), .ZN(
        REG3_1_n53) );
  NAND2_X1 REG3_1_U22 ( .A1(temp3[7]), .A2(REG3_1_n43), .ZN(REG3_1_n82) );
  OAI21_X1 REG3_1_U21 ( .B1(REG3_1_n44), .B2(REG3_1_n69), .A(REG3_1_n82), .ZN(
        REG3_1_n54) );
  NAND2_X1 REG3_1_U20 ( .A1(temp3[6]), .A2(REG3_1_n43), .ZN(REG3_1_n83) );
  OAI21_X1 REG3_1_U19 ( .B1(REG3_1_n44), .B2(REG3_1_n68), .A(REG3_1_n83), .ZN(
        REG3_1_n55) );
  NAND2_X1 REG3_1_U18 ( .A1(temp3[1]), .A2(REG3_1_n43), .ZN(REG3_1_n88) );
  OAI21_X1 REG3_1_U17 ( .B1(REG3_1_n44), .B2(REG3_1_n63), .A(REG3_1_n88), .ZN(
        REG3_1_n60) );
  NAND2_X1 REG3_1_U16 ( .A1(temp3[0]), .A2(REG3_1_n43), .ZN(REG3_1_n89) );
  OAI21_X1 REG3_1_U15 ( .B1(REG3_1_n44), .B2(REG3_1_n62), .A(REG3_1_n89), .ZN(
        REG3_1_n61) );
  NAND2_X1 REG3_1_U14 ( .A1(temp3[10]), .A2(REG3_1_n44), .ZN(REG3_1_n79) );
  OAI21_X1 REG3_1_U13 ( .B1(REG3_1_n44), .B2(REG3_1_n72), .A(REG3_1_n79), .ZN(
        REG3_1_n51) );
  NAND2_X1 REG3_1_U12 ( .A1(temp3[12]), .A2(REG3_1_n43), .ZN(REG3_1_n77) );
  OAI21_X1 REG3_1_U11 ( .B1(REG3_1_n44), .B2(REG3_1_n74), .A(REG3_1_n77), .ZN(
        REG3_1_n49) );
  NAND2_X1 REG3_1_U10 ( .A1(temp3[11]), .A2(REG3_1_n43), .ZN(REG3_1_n78) );
  OAI21_X1 REG3_1_U9 ( .B1(REG3_1_n44), .B2(REG3_1_n73), .A(REG3_1_n78), .ZN(
        REG3_1_n50) );
  NAND2_X1 REG3_1_U8 ( .A1(temp3[13]), .A2(REG3_1_n43), .ZN(REG3_1_n76) );
  OAI21_X1 REG3_1_U7 ( .B1(REG3_1_n44), .B2(REG3_1_n75), .A(REG3_1_n76), .ZN(
        REG3_1_n48) );
  BUF_X1 REG3_1_U6 ( .A(n47), .Z(REG3_1_n47) );
  BUF_X1 REG3_1_U5 ( .A(n47), .Z(REG3_1_n46) );
  BUF_X1 REG3_1_U4 ( .A(VIN), .Z(REG3_1_n45) );
  BUF_X1 REG3_1_U3 ( .A(VIN), .Z(REG3_1_n43) );
  BUF_X1 REG3_1_U2 ( .A(VIN), .Z(REG3_1_n44) );
  DFFR_X1 REG3_1_q_reg_0_ ( .D(REG3_1_n61), .CK(CLK), .RN(REG3_1_n47), .Q(
        mul3_reg[0]), .QN(REG3_1_n62) );
  DFFR_X1 REG3_1_q_reg_1_ ( .D(REG3_1_n60), .CK(CLK), .RN(REG3_1_n47), .Q(
        mul3_reg[1]), .QN(REG3_1_n63) );
  DFFR_X1 REG3_1_q_reg_2_ ( .D(REG3_1_n59), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[2]), .QN(REG3_1_n64) );
  DFFR_X1 REG3_1_q_reg_3_ ( .D(REG3_1_n58), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[3]), .QN(REG3_1_n65) );
  DFFR_X1 REG3_1_q_reg_4_ ( .D(REG3_1_n57), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[4]), .QN(REG3_1_n66) );
  DFFR_X1 REG3_1_q_reg_5_ ( .D(REG3_1_n56), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[5]), .QN(REG3_1_n67) );
  DFFR_X1 REG3_1_q_reg_6_ ( .D(REG3_1_n55), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[6]), .QN(REG3_1_n68) );
  DFFR_X1 REG3_1_q_reg_7_ ( .D(REG3_1_n54), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[7]), .QN(REG3_1_n69) );
  DFFR_X1 REG3_1_q_reg_8_ ( .D(REG3_1_n53), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[8]), .QN(REG3_1_n70) );
  DFFR_X1 REG3_1_q_reg_9_ ( .D(REG3_1_n52), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[9]), .QN(REG3_1_n71) );
  DFFR_X1 REG3_1_q_reg_10_ ( .D(REG3_1_n51), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[10]), .QN(REG3_1_n72) );
  DFFR_X1 REG3_1_q_reg_11_ ( .D(REG3_1_n50), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[11]), .QN(REG3_1_n73) );
  DFFR_X1 REG3_1_q_reg_12_ ( .D(REG3_1_n49), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[12]), .QN(REG3_1_n74) );
  DFFR_X1 REG3_1_q_reg_13_ ( .D(REG3_1_n48), .CK(CLK), .RN(REG3_1_n46), .Q(
        mul3_reg[13]), .QN(REG3_1_n75) );
  NAND2_X1 REGISTER4_U34 ( .A1(reg5[13]), .A2(REGISTER4_n43), .ZN(
        REGISTER4_n76) );
  OAI21_X1 REGISTER4_U33 ( .B1(REGISTER4_n44), .B2(REGISTER4_n75), .A(
        REGISTER4_n76), .ZN(REGISTER4_n48) );
  NAND2_X1 REGISTER4_U32 ( .A1(reg5[12]), .A2(REGISTER4_n43), .ZN(
        REGISTER4_n77) );
  OAI21_X1 REGISTER4_U31 ( .B1(REGISTER4_n44), .B2(REGISTER4_n74), .A(
        REGISTER4_n77), .ZN(REGISTER4_n49) );
  NAND2_X1 REGISTER4_U30 ( .A1(reg5[11]), .A2(REGISTER4_n43), .ZN(
        REGISTER4_n78) );
  OAI21_X1 REGISTER4_U29 ( .B1(REGISTER4_n44), .B2(REGISTER4_n73), .A(
        REGISTER4_n78), .ZN(REGISTER4_n50) );
  NAND2_X1 REGISTER4_U28 ( .A1(reg5[9]), .A2(REGISTER4_n43), .ZN(REGISTER4_n80) );
  OAI21_X1 REGISTER4_U27 ( .B1(REGISTER4_n44), .B2(REGISTER4_n71), .A(
        REGISTER4_n80), .ZN(REGISTER4_n52) );
  NAND2_X1 REGISTER4_U26 ( .A1(reg5[7]), .A2(REGISTER4_n43), .ZN(REGISTER4_n82) );
  OAI21_X1 REGISTER4_U25 ( .B1(REGISTER4_n44), .B2(REGISTER4_n69), .A(
        REGISTER4_n82), .ZN(REGISTER4_n54) );
  NAND2_X1 REGISTER4_U24 ( .A1(reg5[6]), .A2(REGISTER4_n43), .ZN(REGISTER4_n83) );
  OAI21_X1 REGISTER4_U23 ( .B1(REGISTER4_n44), .B2(REGISTER4_n68), .A(
        REGISTER4_n83), .ZN(REGISTER4_n55) );
  NAND2_X1 REGISTER4_U22 ( .A1(reg5[5]), .A2(REGISTER4_n43), .ZN(REGISTER4_n84) );
  OAI21_X1 REGISTER4_U21 ( .B1(REGISTER4_n44), .B2(REGISTER4_n67), .A(
        REGISTER4_n84), .ZN(REGISTER4_n56) );
  NAND2_X1 REGISTER4_U20 ( .A1(reg5[4]), .A2(REGISTER4_n43), .ZN(REGISTER4_n85) );
  OAI21_X1 REGISTER4_U19 ( .B1(REGISTER4_n45), .B2(REGISTER4_n66), .A(
        REGISTER4_n85), .ZN(REGISTER4_n57) );
  NAND2_X1 REGISTER4_U18 ( .A1(reg5[3]), .A2(REGISTER4_n43), .ZN(REGISTER4_n86) );
  OAI21_X1 REGISTER4_U17 ( .B1(REGISTER4_n45), .B2(REGISTER4_n65), .A(
        REGISTER4_n86), .ZN(REGISTER4_n58) );
  NAND2_X1 REGISTER4_U16 ( .A1(reg5[2]), .A2(REGISTER4_n43), .ZN(REGISTER4_n87) );
  OAI21_X1 REGISTER4_U15 ( .B1(REGISTER4_n45), .B2(REGISTER4_n64), .A(
        REGISTER4_n87), .ZN(REGISTER4_n59) );
  NAND2_X1 REGISTER4_U14 ( .A1(reg5[1]), .A2(REGISTER4_n43), .ZN(REGISTER4_n88) );
  OAI21_X1 REGISTER4_U13 ( .B1(REGISTER4_n44), .B2(REGISTER4_n63), .A(
        REGISTER4_n88), .ZN(REGISTER4_n60) );
  NAND2_X1 REGISTER4_U12 ( .A1(reg5[0]), .A2(REGISTER4_n43), .ZN(REGISTER4_n89) );
  OAI21_X1 REGISTER4_U11 ( .B1(REGISTER4_n44), .B2(REGISTER4_n62), .A(
        REGISTER4_n89), .ZN(REGISTER4_n61) );
  NAND2_X1 REGISTER4_U10 ( .A1(reg5[10]), .A2(REGISTER4_n44), .ZN(
        REGISTER4_n79) );
  OAI21_X1 REGISTER4_U9 ( .B1(REGISTER4_n44), .B2(REGISTER4_n72), .A(
        REGISTER4_n79), .ZN(REGISTER4_n51) );
  NAND2_X1 REGISTER4_U8 ( .A1(reg5[8]), .A2(REGISTER4_n44), .ZN(REGISTER4_n81)
         );
  OAI21_X1 REGISTER4_U7 ( .B1(REGISTER4_n44), .B2(REGISTER4_n70), .A(
        REGISTER4_n81), .ZN(REGISTER4_n53) );
  BUF_X1 REGISTER4_U6 ( .A(n47), .Z(REGISTER4_n47) );
  BUF_X1 REGISTER4_U5 ( .A(n47), .Z(REGISTER4_n46) );
  BUF_X1 REGISTER4_U4 ( .A(VIN), .Z(REGISTER4_n45) );
  BUF_X1 REGISTER4_U3 ( .A(VIN), .Z(REGISTER4_n43) );
  BUF_X1 REGISTER4_U2 ( .A(VIN), .Z(REGISTER4_n44) );
  DFFR_X1 REGISTER4_q_reg_0_ ( .D(REGISTER4_n61), .CK(CLK), .RN(REGISTER4_n47), 
        .Q(reg4_reg[0]), .QN(REGISTER4_n62) );
  DFFR_X1 REGISTER4_q_reg_1_ ( .D(REGISTER4_n60), .CK(CLK), .RN(REGISTER4_n47), 
        .Q(reg4_reg[1]), .QN(REGISTER4_n63) );
  DFFR_X1 REGISTER4_q_reg_2_ ( .D(REGISTER4_n59), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[2]), .QN(REGISTER4_n64) );
  DFFR_X1 REGISTER4_q_reg_3_ ( .D(REGISTER4_n58), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[3]), .QN(REGISTER4_n65) );
  DFFR_X1 REGISTER4_q_reg_4_ ( .D(REGISTER4_n57), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[4]), .QN(REGISTER4_n66) );
  DFFR_X1 REGISTER4_q_reg_5_ ( .D(REGISTER4_n56), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[5]), .QN(REGISTER4_n67) );
  DFFR_X1 REGISTER4_q_reg_6_ ( .D(REGISTER4_n55), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[6]), .QN(REGISTER4_n68) );
  DFFR_X1 REGISTER4_q_reg_7_ ( .D(REGISTER4_n54), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[7]), .QN(REGISTER4_n69) );
  DFFR_X1 REGISTER4_q_reg_8_ ( .D(REGISTER4_n53), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[8]), .QN(REGISTER4_n70) );
  DFFR_X1 REGISTER4_q_reg_9_ ( .D(REGISTER4_n52), .CK(CLK), .RN(REGISTER4_n46), 
        .Q(reg4_reg[9]), .QN(REGISTER4_n71) );
  DFFR_X1 REGISTER4_q_reg_10_ ( .D(REGISTER4_n51), .CK(CLK), .RN(REGISTER4_n46), .Q(reg4_reg[10]), .QN(REGISTER4_n72) );
  DFFR_X1 REGISTER4_q_reg_11_ ( .D(REGISTER4_n50), .CK(CLK), .RN(REGISTER4_n46), .Q(reg4_reg[11]), .QN(REGISTER4_n73) );
  DFFR_X1 REGISTER4_q_reg_12_ ( .D(REGISTER4_n49), .CK(CLK), .RN(REGISTER4_n46), .Q(reg4_reg[12]), .QN(REGISTER4_n74) );
  DFFR_X1 REGISTER4_q_reg_13_ ( .D(REGISTER4_n48), .CK(CLK), .RN(REGISTER4_n46), .Q(reg4_reg[13]), .QN(REGISTER4_n75) );
  XOR2_X1 p9_mult_21_U691 ( .A(reg4_reg[2]), .B(reg4_reg[1]), .Z(
        p9_mult_21_n798) );
  INV_X1 p9_mult_21_U690 ( .A(reg4_reg[1]), .ZN(p9_mult_21_n655) );
  NOR2_X1 p9_mult_21_U689 ( .A1(p9_mult_21_n655), .A2(B3[1]), .ZN(
        p9_mult_21_n803) );
  INV_X1 p9_mult_21_U688 ( .A(p9_mult_21_n803), .ZN(p9_mult_21_n805) );
  NAND2_X1 p9_mult_21_U687 ( .A1(reg4_reg[1]), .A2(p9_mult_21_n643), .ZN(
        p9_mult_21_n641) );
  XNOR2_X1 p9_mult_21_U686 ( .A(B3[2]), .B(reg4_reg[1]), .ZN(p9_mult_21_n640)
         );
  OAI22_X1 p9_mult_21_U685 ( .A1(p9_mult_21_n805), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n640), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n804) );
  NAND2_X1 p9_mult_21_U684 ( .A1(p9_mult_21_n798), .A2(p9_mult_21_n804), .ZN(
        p9_mult_21_n801) );
  NAND2_X1 p9_mult_21_U683 ( .A1(p9_mult_21_n803), .A2(p9_mult_21_n804), .ZN(
        p9_mult_21_n802) );
  INV_X1 p9_mult_21_U682 ( .A(B3[0]), .ZN(p9_mult_21_n673) );
  MUX2_X1 p9_mult_21_U681 ( .A(p9_mult_21_n801), .B(p9_mult_21_n802), .S(
        p9_mult_21_n673), .Z(p9_mult_21_n800) );
  INV_X1 p9_mult_21_U680 ( .A(p9_mult_21_n800), .ZN(p9_mult_21_n795) );
  INV_X1 p9_mult_21_U679 ( .A(reg4_reg[3]), .ZN(p9_mult_21_n771) );
  XNOR2_X1 p9_mult_21_U678 ( .A(p9_mult_21_n771), .B(reg4_reg[2]), .ZN(
        p9_mult_21_n799) );
  NAND2_X1 p9_mult_21_U677 ( .A1(p9_mult_21_n658), .A2(p9_mult_21_n799), .ZN(
        p9_mult_21_n657) );
  NAND3_X1 p9_mult_21_U676 ( .A1(p9_mult_21_n798), .A2(p9_mult_21_n673), .A3(
        reg4_reg[3]), .ZN(p9_mult_21_n797) );
  OAI21_X1 p9_mult_21_U675 ( .B1(p9_mult_21_n771), .B2(p9_mult_21_n657), .A(
        p9_mult_21_n797), .ZN(p9_mult_21_n796) );
  AOI222_X1 p9_mult_21_U674 ( .A1(p9_mult_21_n795), .A2(p9_mult_21_n316), .B1(
        p9_mult_21_n796), .B2(p9_mult_21_n795), .C1(p9_mult_21_n796), .C2(
        p9_mult_21_n316), .ZN(p9_mult_21_n794) );
  INV_X1 p9_mult_21_U673 ( .A(p9_mult_21_n794), .ZN(p9_mult_21_n793) );
  AOI222_X1 p9_mult_21_U672 ( .A1(p9_mult_21_n793), .A2(p9_mult_21_n314), .B1(
        p9_mult_21_n793), .B2(p9_mult_21_n315), .C1(p9_mult_21_n315), .C2(
        p9_mult_21_n314), .ZN(p9_mult_21_n792) );
  INV_X1 p9_mult_21_U671 ( .A(p9_mult_21_n792), .ZN(p9_mult_21_n791) );
  AOI222_X1 p9_mult_21_U670 ( .A1(p9_mult_21_n791), .A2(p9_mult_21_n310), .B1(
        p9_mult_21_n791), .B2(p9_mult_21_n313), .C1(p9_mult_21_n313), .C2(
        p9_mult_21_n310), .ZN(p9_mult_21_n790) );
  INV_X1 p9_mult_21_U669 ( .A(p9_mult_21_n790), .ZN(p9_mult_21_n789) );
  AOI222_X1 p9_mult_21_U668 ( .A1(p9_mult_21_n789), .A2(p9_mult_21_n306), .B1(
        p9_mult_21_n789), .B2(p9_mult_21_n309), .C1(p9_mult_21_n309), .C2(
        p9_mult_21_n306), .ZN(p9_mult_21_n788) );
  INV_X1 p9_mult_21_U667 ( .A(p9_mult_21_n788), .ZN(p9_mult_21_n787) );
  AOI222_X1 p9_mult_21_U666 ( .A1(p9_mult_21_n787), .A2(p9_mult_21_n300), .B1(
        p9_mult_21_n787), .B2(p9_mult_21_n305), .C1(p9_mult_21_n305), .C2(
        p9_mult_21_n300), .ZN(p9_mult_21_n786) );
  INV_X1 p9_mult_21_U665 ( .A(p9_mult_21_n786), .ZN(p9_mult_21_n785) );
  AOI222_X1 p9_mult_21_U664 ( .A1(p9_mult_21_n785), .A2(p9_mult_21_n294), .B1(
        p9_mult_21_n785), .B2(p9_mult_21_n299), .C1(p9_mult_21_n299), .C2(
        p9_mult_21_n294), .ZN(p9_mult_21_n784) );
  INV_X1 p9_mult_21_U663 ( .A(p9_mult_21_n784), .ZN(p9_mult_21_n783) );
  AOI222_X1 p9_mult_21_U662 ( .A1(p9_mult_21_n783), .A2(p9_mult_21_n286), .B1(
        p9_mult_21_n783), .B2(p9_mult_21_n293), .C1(p9_mult_21_n293), .C2(
        p9_mult_21_n286), .ZN(p9_mult_21_n780) );
  INV_X1 p9_mult_21_U661 ( .A(p9_mult_21_n278), .ZN(p9_mult_21_n781) );
  INV_X1 p9_mult_21_U660 ( .A(p9_mult_21_n285), .ZN(p9_mult_21_n782) );
  OAI222_X1 p9_mult_21_U659 ( .A1(p9_mult_21_n780), .A2(p9_mult_21_n781), .B1(
        p9_mult_21_n780), .B2(p9_mult_21_n782), .C1(p9_mult_21_n782), .C2(
        p9_mult_21_n781), .ZN(p9_mult_21_n779) );
  AOI222_X1 p9_mult_21_U658 ( .A1(p9_mult_21_n779), .A2(p9_mult_21_n268), .B1(
        p9_mult_21_n779), .B2(p9_mult_21_n277), .C1(p9_mult_21_n277), .C2(
        p9_mult_21_n268), .ZN(p9_mult_21_n776) );
  INV_X1 p9_mult_21_U657 ( .A(p9_mult_21_n258), .ZN(p9_mult_21_n777) );
  INV_X1 p9_mult_21_U656 ( .A(p9_mult_21_n267), .ZN(p9_mult_21_n778) );
  OAI222_X1 p9_mult_21_U655 ( .A1(p9_mult_21_n776), .A2(p9_mult_21_n777), .B1(
        p9_mult_21_n776), .B2(p9_mult_21_n778), .C1(p9_mult_21_n778), .C2(
        p9_mult_21_n777), .ZN(p9_mult_21_n149) );
  XOR2_X1 p9_mult_21_U654 ( .A(B3[12]), .B(reg4_reg[13]), .Z(p9_mult_21_n757)
         );
  INV_X1 p9_mult_21_U653 ( .A(reg4_reg[11]), .ZN(p9_mult_21_n764) );
  INV_X1 p9_mult_21_U652 ( .A(reg4_reg[13]), .ZN(p9_mult_21_n766) );
  XNOR2_X1 p9_mult_21_U651 ( .A(p9_mult_21_n766), .B(reg4_reg[12]), .ZN(
        p9_mult_21_n775) );
  NAND2_X1 p9_mult_21_U650 ( .A1(p9_mult_21_n742), .A2(p9_mult_21_n775), .ZN(
        p9_mult_21_n744) );
  INV_X1 p9_mult_21_U649 ( .A(p9_mult_21_n744), .ZN(p9_mult_21_n637) );
  INV_X1 p9_mult_21_U648 ( .A(p9_mult_21_n742), .ZN(p9_mult_21_n638) );
  XNOR2_X1 p9_mult_21_U647 ( .A(B3[13]), .B(p9_mult_21_n766), .ZN(
        p9_mult_21_n639) );
  AOI22_X1 p9_mult_21_U646 ( .A1(p9_mult_21_n757), .A2(p9_mult_21_n637), .B1(
        p9_mult_21_n638), .B2(p9_mult_21_n639), .ZN(p9_mult_21_n162) );
  XNOR2_X1 p9_mult_21_U645 ( .A(B3[12]), .B(reg4_reg[11]), .ZN(p9_mult_21_n739) );
  INV_X1 p9_mult_21_U644 ( .A(reg4_reg[9]), .ZN(p9_mult_21_n762) );
  XNOR2_X1 p9_mult_21_U643 ( .A(p9_mult_21_n764), .B(reg4_reg[10]), .ZN(
        p9_mult_21_n774) );
  NAND2_X1 p9_mult_21_U642 ( .A1(p9_mult_21_n725), .A2(p9_mult_21_n774), .ZN(
        p9_mult_21_n727) );
  XNOR2_X1 p9_mult_21_U641 ( .A(B3[13]), .B(reg4_reg[11]), .ZN(p9_mult_21_n741) );
  OAI22_X1 p9_mult_21_U640 ( .A1(p9_mult_21_n739), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n741), .ZN(p9_mult_21_n167) );
  INV_X1 p9_mult_21_U639 ( .A(p9_mult_21_n167), .ZN(p9_mult_21_n168) );
  XNOR2_X1 p9_mult_21_U638 ( .A(B3[12]), .B(reg4_reg[9]), .ZN(p9_mult_21_n722)
         );
  INV_X1 p9_mult_21_U637 ( .A(reg4_reg[7]), .ZN(p9_mult_21_n760) );
  XNOR2_X1 p9_mult_21_U636 ( .A(p9_mult_21_n762), .B(reg4_reg[8]), .ZN(
        p9_mult_21_n773) );
  NAND2_X1 p9_mult_21_U635 ( .A1(p9_mult_21_n708), .A2(p9_mult_21_n773), .ZN(
        p9_mult_21_n710) );
  XNOR2_X1 p9_mult_21_U634 ( .A(B3[13]), .B(reg4_reg[9]), .ZN(p9_mult_21_n724)
         );
  OAI22_X1 p9_mult_21_U633 ( .A1(p9_mult_21_n722), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n724), .ZN(p9_mult_21_n177) );
  INV_X1 p9_mult_21_U632 ( .A(p9_mult_21_n177), .ZN(p9_mult_21_n178) );
  XNOR2_X1 p9_mult_21_U631 ( .A(B3[12]), .B(reg4_reg[7]), .ZN(p9_mult_21_n705)
         );
  INV_X1 p9_mult_21_U630 ( .A(reg4_reg[5]), .ZN(p9_mult_21_n758) );
  XNOR2_X1 p9_mult_21_U629 ( .A(p9_mult_21_n760), .B(reg4_reg[6]), .ZN(
        p9_mult_21_n772) );
  NAND2_X1 p9_mult_21_U628 ( .A1(p9_mult_21_n691), .A2(p9_mult_21_n772), .ZN(
        p9_mult_21_n693) );
  XNOR2_X1 p9_mult_21_U627 ( .A(B3[13]), .B(reg4_reg[7]), .ZN(p9_mult_21_n707)
         );
  OAI22_X1 p9_mult_21_U626 ( .A1(p9_mult_21_n705), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n707), .ZN(p9_mult_21_n191) );
  INV_X1 p9_mult_21_U625 ( .A(p9_mult_21_n191), .ZN(p9_mult_21_n192) );
  XNOR2_X1 p9_mult_21_U624 ( .A(B3[12]), .B(reg4_reg[5]), .ZN(p9_mult_21_n688)
         );
  XNOR2_X1 p9_mult_21_U623 ( .A(p9_mult_21_n758), .B(reg4_reg[4]), .ZN(
        p9_mult_21_n770) );
  NAND2_X1 p9_mult_21_U622 ( .A1(p9_mult_21_n674), .A2(p9_mult_21_n770), .ZN(
        p9_mult_21_n676) );
  XNOR2_X1 p9_mult_21_U621 ( .A(B3[13]), .B(reg4_reg[5]), .ZN(p9_mult_21_n690)
         );
  OAI22_X1 p9_mult_21_U620 ( .A1(p9_mult_21_n688), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n690), .ZN(p9_mult_21_n209) );
  INV_X1 p9_mult_21_U619 ( .A(p9_mult_21_n209), .ZN(p9_mult_21_n210) );
  XNOR2_X1 p9_mult_21_U618 ( .A(B3[12]), .B(reg4_reg[3]), .ZN(p9_mult_21_n670)
         );
  XNOR2_X1 p9_mult_21_U617 ( .A(B3[13]), .B(reg4_reg[3]), .ZN(p9_mult_21_n672)
         );
  OAI22_X1 p9_mult_21_U616 ( .A1(p9_mult_21_n670), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n672), .ZN(p9_mult_21_n231) );
  INV_X1 p9_mult_21_U615 ( .A(p9_mult_21_n231), .ZN(p9_mult_21_n232) );
  XNOR2_X1 p9_mult_21_U614 ( .A(B3[3]), .B(reg4_reg[11]), .ZN(p9_mult_21_n730)
         );
  XNOR2_X1 p9_mult_21_U613 ( .A(B3[4]), .B(reg4_reg[11]), .ZN(p9_mult_21_n731)
         );
  OAI22_X1 p9_mult_21_U612 ( .A1(p9_mult_21_n730), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n731), .ZN(p9_mult_21_n768) );
  XNOR2_X1 p9_mult_21_U611 ( .A(B3[9]), .B(reg4_reg[5]), .ZN(p9_mult_21_n685)
         );
  XNOR2_X1 p9_mult_21_U610 ( .A(B3[10]), .B(reg4_reg[5]), .ZN(p9_mult_21_n686)
         );
  OAI22_X1 p9_mult_21_U609 ( .A1(p9_mult_21_n685), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n686), .ZN(p9_mult_21_n769) );
  OR2_X1 p9_mult_21_U608 ( .A1(p9_mult_21_n768), .A2(p9_mult_21_n769), .ZN(
        p9_mult_21_n243) );
  XNOR2_X1 p9_mult_21_U607 ( .A(p9_mult_21_n768), .B(p9_mult_21_n769), .ZN(
        p9_mult_21_n244) );
  NAND3_X1 p9_mult_21_U606 ( .A1(p9_mult_21_n638), .A2(p9_mult_21_n673), .A3(
        reg4_reg[13]), .ZN(p9_mult_21_n767) );
  OAI21_X1 p9_mult_21_U605 ( .B1(p9_mult_21_n766), .B2(p9_mult_21_n744), .A(
        p9_mult_21_n767), .ZN(p9_mult_21_n317) );
  OR3_X1 p9_mult_21_U604 ( .A1(p9_mult_21_n725), .A2(B3[0]), .A3(
        p9_mult_21_n764), .ZN(p9_mult_21_n765) );
  OAI21_X1 p9_mult_21_U603 ( .B1(p9_mult_21_n764), .B2(p9_mult_21_n727), .A(
        p9_mult_21_n765), .ZN(p9_mult_21_n318) );
  OR3_X1 p9_mult_21_U602 ( .A1(p9_mult_21_n708), .A2(B3[0]), .A3(
        p9_mult_21_n762), .ZN(p9_mult_21_n763) );
  OAI21_X1 p9_mult_21_U601 ( .B1(p9_mult_21_n762), .B2(p9_mult_21_n710), .A(
        p9_mult_21_n763), .ZN(p9_mult_21_n319) );
  OR3_X1 p9_mult_21_U600 ( .A1(p9_mult_21_n691), .A2(B3[0]), .A3(
        p9_mult_21_n760), .ZN(p9_mult_21_n761) );
  OAI21_X1 p9_mult_21_U599 ( .B1(p9_mult_21_n760), .B2(p9_mult_21_n693), .A(
        p9_mult_21_n761), .ZN(p9_mult_21_n320) );
  OR3_X1 p9_mult_21_U598 ( .A1(p9_mult_21_n674), .A2(B3[0]), .A3(
        p9_mult_21_n758), .ZN(p9_mult_21_n759) );
  OAI21_X1 p9_mult_21_U597 ( .B1(p9_mult_21_n758), .B2(p9_mult_21_n676), .A(
        p9_mult_21_n759), .ZN(p9_mult_21_n321) );
  XNOR2_X1 p9_mult_21_U596 ( .A(B3[11]), .B(reg4_reg[13]), .ZN(p9_mult_21_n755) );
  INV_X1 p9_mult_21_U595 ( .A(p9_mult_21_n757), .ZN(p9_mult_21_n756) );
  OAI22_X1 p9_mult_21_U594 ( .A1(p9_mult_21_n755), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n756), .ZN(p9_mult_21_n325) );
  XNOR2_X1 p9_mult_21_U593 ( .A(B3[10]), .B(reg4_reg[13]), .ZN(p9_mult_21_n754) );
  OAI22_X1 p9_mult_21_U592 ( .A1(p9_mult_21_n754), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n755), .ZN(p9_mult_21_n326) );
  XNOR2_X1 p9_mult_21_U591 ( .A(B3[9]), .B(reg4_reg[13]), .ZN(p9_mult_21_n753)
         );
  OAI22_X1 p9_mult_21_U590 ( .A1(p9_mult_21_n753), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n754), .ZN(p9_mult_21_n327) );
  XNOR2_X1 p9_mult_21_U589 ( .A(B3[8]), .B(reg4_reg[13]), .ZN(p9_mult_21_n752)
         );
  OAI22_X1 p9_mult_21_U588 ( .A1(p9_mult_21_n752), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n753), .ZN(p9_mult_21_n328) );
  XNOR2_X1 p9_mult_21_U587 ( .A(B3[7]), .B(reg4_reg[13]), .ZN(p9_mult_21_n751)
         );
  OAI22_X1 p9_mult_21_U586 ( .A1(p9_mult_21_n751), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n752), .ZN(p9_mult_21_n329) );
  XNOR2_X1 p9_mult_21_U585 ( .A(B3[6]), .B(reg4_reg[13]), .ZN(p9_mult_21_n750)
         );
  OAI22_X1 p9_mult_21_U584 ( .A1(p9_mult_21_n750), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n751), .ZN(p9_mult_21_n330) );
  XNOR2_X1 p9_mult_21_U583 ( .A(B3[5]), .B(reg4_reg[13]), .ZN(p9_mult_21_n749)
         );
  OAI22_X1 p9_mult_21_U582 ( .A1(p9_mult_21_n749), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n750), .ZN(p9_mult_21_n331) );
  XNOR2_X1 p9_mult_21_U581 ( .A(B3[4]), .B(reg4_reg[13]), .ZN(p9_mult_21_n748)
         );
  OAI22_X1 p9_mult_21_U580 ( .A1(p9_mult_21_n748), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n749), .ZN(p9_mult_21_n332) );
  XNOR2_X1 p9_mult_21_U579 ( .A(B3[3]), .B(reg4_reg[13]), .ZN(p9_mult_21_n747)
         );
  OAI22_X1 p9_mult_21_U578 ( .A1(p9_mult_21_n747), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n748), .ZN(p9_mult_21_n333) );
  XNOR2_X1 p9_mult_21_U577 ( .A(B3[2]), .B(reg4_reg[13]), .ZN(p9_mult_21_n746)
         );
  OAI22_X1 p9_mult_21_U576 ( .A1(p9_mult_21_n746), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n747), .ZN(p9_mult_21_n334) );
  XNOR2_X1 p9_mult_21_U575 ( .A(B3[1]), .B(reg4_reg[13]), .ZN(p9_mult_21_n745)
         );
  OAI22_X1 p9_mult_21_U574 ( .A1(p9_mult_21_n745), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n746), .ZN(p9_mult_21_n335) );
  XNOR2_X1 p9_mult_21_U573 ( .A(reg4_reg[13]), .B(B3[0]), .ZN(p9_mult_21_n743)
         );
  OAI22_X1 p9_mult_21_U572 ( .A1(p9_mult_21_n743), .A2(p9_mult_21_n744), .B1(
        p9_mult_21_n742), .B2(p9_mult_21_n745), .ZN(p9_mult_21_n336) );
  NOR2_X1 p9_mult_21_U571 ( .A1(p9_mult_21_n673), .A2(p9_mult_21_n742), .ZN(
        p9_mult_21_n337) );
  AOI21_X1 p9_mult_21_U570 ( .B1(p9_mult_21_n727), .B2(p9_mult_21_n725), .A(
        p9_mult_21_n741), .ZN(p9_mult_21_n740) );
  INV_X1 p9_mult_21_U569 ( .A(p9_mult_21_n740), .ZN(p9_mult_21_n338) );
  XNOR2_X1 p9_mult_21_U568 ( .A(B3[11]), .B(reg4_reg[11]), .ZN(p9_mult_21_n738) );
  OAI22_X1 p9_mult_21_U567 ( .A1(p9_mult_21_n738), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n739), .ZN(p9_mult_21_n339) );
  XNOR2_X1 p9_mult_21_U566 ( .A(B3[10]), .B(reg4_reg[11]), .ZN(p9_mult_21_n737) );
  OAI22_X1 p9_mult_21_U565 ( .A1(p9_mult_21_n737), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n738), .ZN(p9_mult_21_n340) );
  XNOR2_X1 p9_mult_21_U564 ( .A(B3[9]), .B(reg4_reg[11]), .ZN(p9_mult_21_n736)
         );
  OAI22_X1 p9_mult_21_U563 ( .A1(p9_mult_21_n736), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n737), .ZN(p9_mult_21_n341) );
  XNOR2_X1 p9_mult_21_U562 ( .A(B3[8]), .B(reg4_reg[11]), .ZN(p9_mult_21_n735)
         );
  OAI22_X1 p9_mult_21_U561 ( .A1(p9_mult_21_n735), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n736), .ZN(p9_mult_21_n342) );
  XNOR2_X1 p9_mult_21_U560 ( .A(B3[7]), .B(reg4_reg[11]), .ZN(p9_mult_21_n734)
         );
  OAI22_X1 p9_mult_21_U559 ( .A1(p9_mult_21_n734), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n735), .ZN(p9_mult_21_n343) );
  XNOR2_X1 p9_mult_21_U558 ( .A(B3[6]), .B(reg4_reg[11]), .ZN(p9_mult_21_n733)
         );
  OAI22_X1 p9_mult_21_U557 ( .A1(p9_mult_21_n733), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n734), .ZN(p9_mult_21_n344) );
  XNOR2_X1 p9_mult_21_U556 ( .A(B3[5]), .B(reg4_reg[11]), .ZN(p9_mult_21_n732)
         );
  OAI22_X1 p9_mult_21_U555 ( .A1(p9_mult_21_n732), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n733), .ZN(p9_mult_21_n345) );
  OAI22_X1 p9_mult_21_U554 ( .A1(p9_mult_21_n731), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n732), .ZN(p9_mult_21_n346) );
  XNOR2_X1 p9_mult_21_U553 ( .A(B3[2]), .B(reg4_reg[11]), .ZN(p9_mult_21_n729)
         );
  OAI22_X1 p9_mult_21_U552 ( .A1(p9_mult_21_n729), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n730), .ZN(p9_mult_21_n348) );
  XNOR2_X1 p9_mult_21_U551 ( .A(B3[1]), .B(reg4_reg[11]), .ZN(p9_mult_21_n728)
         );
  OAI22_X1 p9_mult_21_U550 ( .A1(p9_mult_21_n728), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n729), .ZN(p9_mult_21_n349) );
  XNOR2_X1 p9_mult_21_U549 ( .A(reg4_reg[11]), .B(B3[0]), .ZN(p9_mult_21_n726)
         );
  OAI22_X1 p9_mult_21_U548 ( .A1(p9_mult_21_n726), .A2(p9_mult_21_n727), .B1(
        p9_mult_21_n725), .B2(p9_mult_21_n728), .ZN(p9_mult_21_n350) );
  NOR2_X1 p9_mult_21_U547 ( .A1(p9_mult_21_n673), .A2(p9_mult_21_n725), .ZN(
        p9_mult_21_n351) );
  AOI21_X1 p9_mult_21_U546 ( .B1(p9_mult_21_n710), .B2(p9_mult_21_n708), .A(
        p9_mult_21_n724), .ZN(p9_mult_21_n723) );
  INV_X1 p9_mult_21_U545 ( .A(p9_mult_21_n723), .ZN(p9_mult_21_n352) );
  XNOR2_X1 p9_mult_21_U544 ( .A(B3[11]), .B(reg4_reg[9]), .ZN(p9_mult_21_n721)
         );
  OAI22_X1 p9_mult_21_U543 ( .A1(p9_mult_21_n721), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n722), .ZN(p9_mult_21_n353) );
  XNOR2_X1 p9_mult_21_U542 ( .A(B3[10]), .B(reg4_reg[9]), .ZN(p9_mult_21_n720)
         );
  OAI22_X1 p9_mult_21_U541 ( .A1(p9_mult_21_n720), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n721), .ZN(p9_mult_21_n354) );
  XNOR2_X1 p9_mult_21_U540 ( .A(B3[9]), .B(reg4_reg[9]), .ZN(p9_mult_21_n719)
         );
  OAI22_X1 p9_mult_21_U539 ( .A1(p9_mult_21_n719), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n720), .ZN(p9_mult_21_n355) );
  XNOR2_X1 p9_mult_21_U538 ( .A(B3[8]), .B(reg4_reg[9]), .ZN(p9_mult_21_n718)
         );
  OAI22_X1 p9_mult_21_U537 ( .A1(p9_mult_21_n718), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n719), .ZN(p9_mult_21_n356) );
  XNOR2_X1 p9_mult_21_U536 ( .A(B3[7]), .B(reg4_reg[9]), .ZN(p9_mult_21_n717)
         );
  OAI22_X1 p9_mult_21_U535 ( .A1(p9_mult_21_n717), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n718), .ZN(p9_mult_21_n357) );
  XNOR2_X1 p9_mult_21_U534 ( .A(B3[6]), .B(reg4_reg[9]), .ZN(p9_mult_21_n716)
         );
  OAI22_X1 p9_mult_21_U533 ( .A1(p9_mult_21_n716), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n717), .ZN(p9_mult_21_n358) );
  XNOR2_X1 p9_mult_21_U532 ( .A(B3[5]), .B(reg4_reg[9]), .ZN(p9_mult_21_n715)
         );
  OAI22_X1 p9_mult_21_U531 ( .A1(p9_mult_21_n715), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n716), .ZN(p9_mult_21_n359) );
  XNOR2_X1 p9_mult_21_U530 ( .A(B3[4]), .B(reg4_reg[9]), .ZN(p9_mult_21_n714)
         );
  OAI22_X1 p9_mult_21_U529 ( .A1(p9_mult_21_n714), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n715), .ZN(p9_mult_21_n360) );
  XNOR2_X1 p9_mult_21_U528 ( .A(B3[3]), .B(reg4_reg[9]), .ZN(p9_mult_21_n713)
         );
  OAI22_X1 p9_mult_21_U527 ( .A1(p9_mult_21_n713), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n714), .ZN(p9_mult_21_n361) );
  XNOR2_X1 p9_mult_21_U526 ( .A(B3[2]), .B(reg4_reg[9]), .ZN(p9_mult_21_n712)
         );
  OAI22_X1 p9_mult_21_U525 ( .A1(p9_mult_21_n712), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n713), .ZN(p9_mult_21_n362) );
  XNOR2_X1 p9_mult_21_U524 ( .A(B3[1]), .B(reg4_reg[9]), .ZN(p9_mult_21_n711)
         );
  OAI22_X1 p9_mult_21_U523 ( .A1(p9_mult_21_n711), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n712), .ZN(p9_mult_21_n363) );
  XNOR2_X1 p9_mult_21_U522 ( .A(reg4_reg[9]), .B(B3[0]), .ZN(p9_mult_21_n709)
         );
  OAI22_X1 p9_mult_21_U521 ( .A1(p9_mult_21_n709), .A2(p9_mult_21_n710), .B1(
        p9_mult_21_n708), .B2(p9_mult_21_n711), .ZN(p9_mult_21_n364) );
  NOR2_X1 p9_mult_21_U520 ( .A1(p9_mult_21_n673), .A2(p9_mult_21_n708), .ZN(
        p9_mult_21_n365) );
  AOI21_X1 p9_mult_21_U519 ( .B1(p9_mult_21_n693), .B2(p9_mult_21_n691), .A(
        p9_mult_21_n707), .ZN(p9_mult_21_n706) );
  INV_X1 p9_mult_21_U518 ( .A(p9_mult_21_n706), .ZN(p9_mult_21_n366) );
  XNOR2_X1 p9_mult_21_U517 ( .A(B3[11]), .B(reg4_reg[7]), .ZN(p9_mult_21_n704)
         );
  OAI22_X1 p9_mult_21_U516 ( .A1(p9_mult_21_n704), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n705), .ZN(p9_mult_21_n367) );
  XNOR2_X1 p9_mult_21_U515 ( .A(B3[10]), .B(reg4_reg[7]), .ZN(p9_mult_21_n703)
         );
  OAI22_X1 p9_mult_21_U514 ( .A1(p9_mult_21_n703), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n704), .ZN(p9_mult_21_n368) );
  XNOR2_X1 p9_mult_21_U513 ( .A(B3[9]), .B(reg4_reg[7]), .ZN(p9_mult_21_n702)
         );
  OAI22_X1 p9_mult_21_U512 ( .A1(p9_mult_21_n702), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n703), .ZN(p9_mult_21_n369) );
  XNOR2_X1 p9_mult_21_U511 ( .A(B3[8]), .B(reg4_reg[7]), .ZN(p9_mult_21_n701)
         );
  OAI22_X1 p9_mult_21_U510 ( .A1(p9_mult_21_n701), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n702), .ZN(p9_mult_21_n370) );
  XNOR2_X1 p9_mult_21_U509 ( .A(B3[7]), .B(reg4_reg[7]), .ZN(p9_mult_21_n700)
         );
  OAI22_X1 p9_mult_21_U508 ( .A1(p9_mult_21_n700), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n701), .ZN(p9_mult_21_n371) );
  XNOR2_X1 p9_mult_21_U507 ( .A(B3[6]), .B(reg4_reg[7]), .ZN(p9_mult_21_n699)
         );
  OAI22_X1 p9_mult_21_U506 ( .A1(p9_mult_21_n699), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n700), .ZN(p9_mult_21_n372) );
  XNOR2_X1 p9_mult_21_U505 ( .A(B3[5]), .B(reg4_reg[7]), .ZN(p9_mult_21_n698)
         );
  OAI22_X1 p9_mult_21_U504 ( .A1(p9_mult_21_n698), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n699), .ZN(p9_mult_21_n373) );
  XNOR2_X1 p9_mult_21_U503 ( .A(B3[4]), .B(reg4_reg[7]), .ZN(p9_mult_21_n697)
         );
  OAI22_X1 p9_mult_21_U502 ( .A1(p9_mult_21_n697), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n698), .ZN(p9_mult_21_n374) );
  XNOR2_X1 p9_mult_21_U501 ( .A(B3[3]), .B(reg4_reg[7]), .ZN(p9_mult_21_n696)
         );
  OAI22_X1 p9_mult_21_U500 ( .A1(p9_mult_21_n696), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n697), .ZN(p9_mult_21_n375) );
  XNOR2_X1 p9_mult_21_U499 ( .A(B3[2]), .B(reg4_reg[7]), .ZN(p9_mult_21_n695)
         );
  OAI22_X1 p9_mult_21_U498 ( .A1(p9_mult_21_n695), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n696), .ZN(p9_mult_21_n376) );
  XNOR2_X1 p9_mult_21_U497 ( .A(B3[1]), .B(reg4_reg[7]), .ZN(p9_mult_21_n694)
         );
  OAI22_X1 p9_mult_21_U496 ( .A1(p9_mult_21_n694), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n695), .ZN(p9_mult_21_n377) );
  XNOR2_X1 p9_mult_21_U495 ( .A(reg4_reg[7]), .B(B3[0]), .ZN(p9_mult_21_n692)
         );
  OAI22_X1 p9_mult_21_U494 ( .A1(p9_mult_21_n692), .A2(p9_mult_21_n693), .B1(
        p9_mult_21_n691), .B2(p9_mult_21_n694), .ZN(p9_mult_21_n378) );
  NOR2_X1 p9_mult_21_U493 ( .A1(p9_mult_21_n673), .A2(p9_mult_21_n691), .ZN(
        p9_mult_21_n379) );
  AOI21_X1 p9_mult_21_U492 ( .B1(p9_mult_21_n676), .B2(p9_mult_21_n674), .A(
        p9_mult_21_n690), .ZN(p9_mult_21_n689) );
  INV_X1 p9_mult_21_U491 ( .A(p9_mult_21_n689), .ZN(p9_mult_21_n380) );
  XNOR2_X1 p9_mult_21_U490 ( .A(B3[11]), .B(reg4_reg[5]), .ZN(p9_mult_21_n687)
         );
  OAI22_X1 p9_mult_21_U489 ( .A1(p9_mult_21_n687), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n688), .ZN(p9_mult_21_n381) );
  OAI22_X1 p9_mult_21_U488 ( .A1(p9_mult_21_n686), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n687), .ZN(p9_mult_21_n382) );
  XNOR2_X1 p9_mult_21_U487 ( .A(B3[8]), .B(reg4_reg[5]), .ZN(p9_mult_21_n684)
         );
  OAI22_X1 p9_mult_21_U486 ( .A1(p9_mult_21_n684), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n685), .ZN(p9_mult_21_n384) );
  XNOR2_X1 p9_mult_21_U485 ( .A(B3[7]), .B(reg4_reg[5]), .ZN(p9_mult_21_n683)
         );
  OAI22_X1 p9_mult_21_U484 ( .A1(p9_mult_21_n683), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n684), .ZN(p9_mult_21_n385) );
  XNOR2_X1 p9_mult_21_U483 ( .A(B3[6]), .B(reg4_reg[5]), .ZN(p9_mult_21_n682)
         );
  OAI22_X1 p9_mult_21_U482 ( .A1(p9_mult_21_n682), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n683), .ZN(p9_mult_21_n386) );
  XNOR2_X1 p9_mult_21_U481 ( .A(B3[5]), .B(reg4_reg[5]), .ZN(p9_mult_21_n681)
         );
  OAI22_X1 p9_mult_21_U480 ( .A1(p9_mult_21_n681), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n682), .ZN(p9_mult_21_n387) );
  XNOR2_X1 p9_mult_21_U479 ( .A(B3[4]), .B(reg4_reg[5]), .ZN(p9_mult_21_n680)
         );
  OAI22_X1 p9_mult_21_U478 ( .A1(p9_mult_21_n680), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n681), .ZN(p9_mult_21_n388) );
  XNOR2_X1 p9_mult_21_U477 ( .A(B3[3]), .B(reg4_reg[5]), .ZN(p9_mult_21_n679)
         );
  OAI22_X1 p9_mult_21_U476 ( .A1(p9_mult_21_n679), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n680), .ZN(p9_mult_21_n389) );
  XNOR2_X1 p9_mult_21_U475 ( .A(B3[2]), .B(reg4_reg[5]), .ZN(p9_mult_21_n678)
         );
  OAI22_X1 p9_mult_21_U474 ( .A1(p9_mult_21_n678), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n679), .ZN(p9_mult_21_n390) );
  XNOR2_X1 p9_mult_21_U473 ( .A(B3[1]), .B(reg4_reg[5]), .ZN(p9_mult_21_n677)
         );
  OAI22_X1 p9_mult_21_U472 ( .A1(p9_mult_21_n677), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n678), .ZN(p9_mult_21_n391) );
  XNOR2_X1 p9_mult_21_U471 ( .A(reg4_reg[5]), .B(B3[0]), .ZN(p9_mult_21_n675)
         );
  OAI22_X1 p9_mult_21_U470 ( .A1(p9_mult_21_n675), .A2(p9_mult_21_n676), .B1(
        p9_mult_21_n674), .B2(p9_mult_21_n677), .ZN(p9_mult_21_n392) );
  NOR2_X1 p9_mult_21_U469 ( .A1(p9_mult_21_n673), .A2(p9_mult_21_n674), .ZN(
        p9_mult_21_n393) );
  AOI21_X1 p9_mult_21_U468 ( .B1(p9_mult_21_n657), .B2(p9_mult_21_n658), .A(
        p9_mult_21_n672), .ZN(p9_mult_21_n671) );
  INV_X1 p9_mult_21_U467 ( .A(p9_mult_21_n671), .ZN(p9_mult_21_n394) );
  XNOR2_X1 p9_mult_21_U466 ( .A(B3[11]), .B(reg4_reg[3]), .ZN(p9_mult_21_n669)
         );
  OAI22_X1 p9_mult_21_U465 ( .A1(p9_mult_21_n669), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n670), .ZN(p9_mult_21_n395) );
  XNOR2_X1 p9_mult_21_U464 ( .A(B3[10]), .B(reg4_reg[3]), .ZN(p9_mult_21_n668)
         );
  OAI22_X1 p9_mult_21_U463 ( .A1(p9_mult_21_n668), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n669), .ZN(p9_mult_21_n396) );
  XNOR2_X1 p9_mult_21_U462 ( .A(B3[9]), .B(reg4_reg[3]), .ZN(p9_mult_21_n667)
         );
  OAI22_X1 p9_mult_21_U461 ( .A1(p9_mult_21_n667), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n668), .ZN(p9_mult_21_n397) );
  XNOR2_X1 p9_mult_21_U460 ( .A(B3[8]), .B(reg4_reg[3]), .ZN(p9_mult_21_n666)
         );
  OAI22_X1 p9_mult_21_U459 ( .A1(p9_mult_21_n666), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n667), .ZN(p9_mult_21_n398) );
  XNOR2_X1 p9_mult_21_U458 ( .A(B3[7]), .B(reg4_reg[3]), .ZN(p9_mult_21_n665)
         );
  OAI22_X1 p9_mult_21_U457 ( .A1(p9_mult_21_n665), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n666), .ZN(p9_mult_21_n399) );
  XNOR2_X1 p9_mult_21_U456 ( .A(B3[6]), .B(reg4_reg[3]), .ZN(p9_mult_21_n664)
         );
  OAI22_X1 p9_mult_21_U455 ( .A1(p9_mult_21_n664), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n665), .ZN(p9_mult_21_n400) );
  XNOR2_X1 p9_mult_21_U454 ( .A(B3[5]), .B(reg4_reg[3]), .ZN(p9_mult_21_n663)
         );
  OAI22_X1 p9_mult_21_U453 ( .A1(p9_mult_21_n663), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n664), .ZN(p9_mult_21_n401) );
  XNOR2_X1 p9_mult_21_U452 ( .A(B3[4]), .B(reg4_reg[3]), .ZN(p9_mult_21_n662)
         );
  OAI22_X1 p9_mult_21_U451 ( .A1(p9_mult_21_n662), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n663), .ZN(p9_mult_21_n402) );
  XNOR2_X1 p9_mult_21_U450 ( .A(B3[3]), .B(reg4_reg[3]), .ZN(p9_mult_21_n661)
         );
  OAI22_X1 p9_mult_21_U449 ( .A1(p9_mult_21_n661), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n662), .ZN(p9_mult_21_n403) );
  XNOR2_X1 p9_mult_21_U448 ( .A(B3[2]), .B(reg4_reg[3]), .ZN(p9_mult_21_n660)
         );
  OAI22_X1 p9_mult_21_U447 ( .A1(p9_mult_21_n660), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n661), .ZN(p9_mult_21_n404) );
  XNOR2_X1 p9_mult_21_U446 ( .A(B3[1]), .B(reg4_reg[3]), .ZN(p9_mult_21_n659)
         );
  OAI22_X1 p9_mult_21_U445 ( .A1(p9_mult_21_n659), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n660), .ZN(p9_mult_21_n405) );
  XNOR2_X1 p9_mult_21_U444 ( .A(reg4_reg[3]), .B(B3[0]), .ZN(p9_mult_21_n656)
         );
  OAI22_X1 p9_mult_21_U443 ( .A1(p9_mult_21_n656), .A2(p9_mult_21_n657), .B1(
        p9_mult_21_n658), .B2(p9_mult_21_n659), .ZN(p9_mult_21_n406) );
  XOR2_X1 p9_mult_21_U442 ( .A(B3[13]), .B(p9_mult_21_n655), .Z(
        p9_mult_21_n653) );
  AOI21_X1 p9_mult_21_U441 ( .B1(p9_mult_21_n641), .B2(p9_mult_21_n643), .A(
        p9_mult_21_n653), .ZN(p9_mult_21_n654) );
  INV_X1 p9_mult_21_U440 ( .A(p9_mult_21_n654), .ZN(p9_mult_21_n408) );
  XNOR2_X1 p9_mult_21_U439 ( .A(B3[12]), .B(reg4_reg[1]), .ZN(p9_mult_21_n652)
         );
  OAI22_X1 p9_mult_21_U438 ( .A1(p9_mult_21_n652), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n653), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n409) );
  XNOR2_X1 p9_mult_21_U437 ( .A(B3[11]), .B(reg4_reg[1]), .ZN(p9_mult_21_n651)
         );
  OAI22_X1 p9_mult_21_U436 ( .A1(p9_mult_21_n651), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n652), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n410) );
  XNOR2_X1 p9_mult_21_U435 ( .A(B3[10]), .B(reg4_reg[1]), .ZN(p9_mult_21_n650)
         );
  OAI22_X1 p9_mult_21_U434 ( .A1(p9_mult_21_n650), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n651), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n411) );
  XNOR2_X1 p9_mult_21_U433 ( .A(B3[9]), .B(reg4_reg[1]), .ZN(p9_mult_21_n649)
         );
  OAI22_X1 p9_mult_21_U432 ( .A1(p9_mult_21_n649), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n650), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n412) );
  XNOR2_X1 p9_mult_21_U431 ( .A(B3[8]), .B(reg4_reg[1]), .ZN(p9_mult_21_n648)
         );
  OAI22_X1 p9_mult_21_U430 ( .A1(p9_mult_21_n648), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n649), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n413) );
  XNOR2_X1 p9_mult_21_U429 ( .A(B3[7]), .B(reg4_reg[1]), .ZN(p9_mult_21_n647)
         );
  OAI22_X1 p9_mult_21_U428 ( .A1(p9_mult_21_n647), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n648), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n414) );
  XNOR2_X1 p9_mult_21_U427 ( .A(B3[6]), .B(reg4_reg[1]), .ZN(p9_mult_21_n646)
         );
  OAI22_X1 p9_mult_21_U426 ( .A1(p9_mult_21_n646), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n647), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n415) );
  XNOR2_X1 p9_mult_21_U425 ( .A(B3[5]), .B(reg4_reg[1]), .ZN(p9_mult_21_n645)
         );
  OAI22_X1 p9_mult_21_U424 ( .A1(p9_mult_21_n645), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n646), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n416) );
  XNOR2_X1 p9_mult_21_U423 ( .A(B3[4]), .B(reg4_reg[1]), .ZN(p9_mult_21_n644)
         );
  OAI22_X1 p9_mult_21_U422 ( .A1(p9_mult_21_n644), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n645), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n417) );
  XNOR2_X1 p9_mult_21_U421 ( .A(B3[3]), .B(reg4_reg[1]), .ZN(p9_mult_21_n642)
         );
  OAI22_X1 p9_mult_21_U420 ( .A1(p9_mult_21_n642), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n644), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n418) );
  OAI22_X1 p9_mult_21_U419 ( .A1(p9_mult_21_n640), .A2(p9_mult_21_n641), .B1(
        p9_mult_21_n642), .B2(p9_mult_21_n643), .ZN(p9_mult_21_n419) );
  OAI21_X1 p9_mult_21_U418 ( .B1(p9_mult_21_n637), .B2(p9_mult_21_n638), .A(
        p9_mult_21_n639), .ZN(p9_mult_21_n636) );
  XOR2_X1 p9_mult_21_U417 ( .A(p9_mult_21_n636), .B(p9_mult_21_n136), .Z(
        p9_mult_21_n635) );
  XNOR2_X1 p9_mult_21_U416 ( .A(p9_mult_21_n162), .B(p9_mult_21_n635), .ZN(
        temp4[13]) );
  XOR2_X2 p9_mult_21_U415 ( .A(reg4_reg[12]), .B(p9_mult_21_n764), .Z(
        p9_mult_21_n742) );
  XOR2_X2 p9_mult_21_U414 ( .A(reg4_reg[10]), .B(p9_mult_21_n762), .Z(
        p9_mult_21_n725) );
  XOR2_X2 p9_mult_21_U413 ( .A(reg4_reg[8]), .B(p9_mult_21_n760), .Z(
        p9_mult_21_n708) );
  XOR2_X2 p9_mult_21_U412 ( .A(reg4_reg[6]), .B(p9_mult_21_n758), .Z(
        p9_mult_21_n691) );
  XOR2_X2 p9_mult_21_U411 ( .A(reg4_reg[4]), .B(p9_mult_21_n771), .Z(
        p9_mult_21_n674) );
  INV_X1 p9_mult_21_U410 ( .A(reg4_reg[0]), .ZN(p9_mult_21_n643) );
  INV_X1 p9_mult_21_U409 ( .A(p9_mult_21_n798), .ZN(p9_mult_21_n658) );
  HA_X1 p9_mult_21_U145 ( .A(p9_mult_21_n406), .B(p9_mult_21_n419), .CO(
        p9_mult_21_n315), .S(p9_mult_21_n316) );
  FA_X1 p9_mult_21_U144 ( .A(p9_mult_21_n418), .B(p9_mult_21_n393), .CI(
        p9_mult_21_n405), .CO(p9_mult_21_n313), .S(p9_mult_21_n314) );
  HA_X1 p9_mult_21_U143 ( .A(p9_mult_21_n321), .B(p9_mult_21_n392), .CO(
        p9_mult_21_n311), .S(p9_mult_21_n312) );
  FA_X1 p9_mult_21_U142 ( .A(p9_mult_21_n404), .B(p9_mult_21_n417), .CI(
        p9_mult_21_n312), .CO(p9_mult_21_n309), .S(p9_mult_21_n310) );
  FA_X1 p9_mult_21_U141 ( .A(p9_mult_21_n416), .B(p9_mult_21_n379), .CI(
        p9_mult_21_n403), .CO(p9_mult_21_n307), .S(p9_mult_21_n308) );
  FA_X1 p9_mult_21_U140 ( .A(p9_mult_21_n311), .B(p9_mult_21_n391), .CI(
        p9_mult_21_n308), .CO(p9_mult_21_n305), .S(p9_mult_21_n306) );
  HA_X1 p9_mult_21_U139 ( .A(p9_mult_21_n320), .B(p9_mult_21_n378), .CO(
        p9_mult_21_n303), .S(p9_mult_21_n304) );
  FA_X1 p9_mult_21_U138 ( .A(p9_mult_21_n390), .B(p9_mult_21_n415), .CI(
        p9_mult_21_n402), .CO(p9_mult_21_n301), .S(p9_mult_21_n302) );
  FA_X1 p9_mult_21_U137 ( .A(p9_mult_21_n307), .B(p9_mult_21_n304), .CI(
        p9_mult_21_n302), .CO(p9_mult_21_n299), .S(p9_mult_21_n300) );
  FA_X1 p9_mult_21_U136 ( .A(p9_mult_21_n389), .B(p9_mult_21_n365), .CI(
        p9_mult_21_n414), .CO(p9_mult_21_n297), .S(p9_mult_21_n298) );
  FA_X1 p9_mult_21_U135 ( .A(p9_mult_21_n377), .B(p9_mult_21_n401), .CI(
        p9_mult_21_n303), .CO(p9_mult_21_n295), .S(p9_mult_21_n296) );
  FA_X1 p9_mult_21_U134 ( .A(p9_mult_21_n298), .B(p9_mult_21_n301), .CI(
        p9_mult_21_n296), .CO(p9_mult_21_n293), .S(p9_mult_21_n294) );
  HA_X1 p9_mult_21_U133 ( .A(p9_mult_21_n319), .B(p9_mult_21_n364), .CO(
        p9_mult_21_n291), .S(p9_mult_21_n292) );
  FA_X1 p9_mult_21_U132 ( .A(p9_mult_21_n376), .B(p9_mult_21_n388), .CI(
        p9_mult_21_n400), .CO(p9_mult_21_n289), .S(p9_mult_21_n290) );
  FA_X1 p9_mult_21_U131 ( .A(p9_mult_21_n292), .B(p9_mult_21_n413), .CI(
        p9_mult_21_n297), .CO(p9_mult_21_n287), .S(p9_mult_21_n288) );
  FA_X1 p9_mult_21_U130 ( .A(p9_mult_21_n290), .B(p9_mult_21_n295), .CI(
        p9_mult_21_n288), .CO(p9_mult_21_n285), .S(p9_mult_21_n286) );
  FA_X1 p9_mult_21_U129 ( .A(p9_mult_21_n375), .B(p9_mult_21_n351), .CI(
        p9_mult_21_n412), .CO(p9_mult_21_n283), .S(p9_mult_21_n284) );
  FA_X1 p9_mult_21_U128 ( .A(p9_mult_21_n363), .B(p9_mult_21_n399), .CI(
        p9_mult_21_n387), .CO(p9_mult_21_n281), .S(p9_mult_21_n282) );
  FA_X1 p9_mult_21_U127 ( .A(p9_mult_21_n289), .B(p9_mult_21_n291), .CI(
        p9_mult_21_n284), .CO(p9_mult_21_n279), .S(p9_mult_21_n280) );
  FA_X1 p9_mult_21_U126 ( .A(p9_mult_21_n287), .B(p9_mult_21_n282), .CI(
        p9_mult_21_n280), .CO(p9_mult_21_n277), .S(p9_mult_21_n278) );
  HA_X1 p9_mult_21_U125 ( .A(p9_mult_21_n318), .B(p9_mult_21_n350), .CO(
        p9_mult_21_n275), .S(p9_mult_21_n276) );
  FA_X1 p9_mult_21_U124 ( .A(p9_mult_21_n362), .B(p9_mult_21_n386), .CI(
        p9_mult_21_n411), .CO(p9_mult_21_n273), .S(p9_mult_21_n274) );
  FA_X1 p9_mult_21_U123 ( .A(p9_mult_21_n374), .B(p9_mult_21_n398), .CI(
        p9_mult_21_n276), .CO(p9_mult_21_n271), .S(p9_mult_21_n272) );
  FA_X1 p9_mult_21_U122 ( .A(p9_mult_21_n281), .B(p9_mult_21_n283), .CI(
        p9_mult_21_n274), .CO(p9_mult_21_n269), .S(p9_mult_21_n270) );
  FA_X1 p9_mult_21_U121 ( .A(p9_mult_21_n279), .B(p9_mult_21_n272), .CI(
        p9_mult_21_n270), .CO(p9_mult_21_n267), .S(p9_mult_21_n268) );
  FA_X1 p9_mult_21_U120 ( .A(p9_mult_21_n361), .B(p9_mult_21_n337), .CI(
        p9_mult_21_n410), .CO(p9_mult_21_n265), .S(p9_mult_21_n266) );
  FA_X1 p9_mult_21_U109 ( .A(p9_mult_21_n349), .B(p9_mult_21_n397), .CI(
        p9_mult_21_n373), .CO(p9_mult_21_n263), .S(p9_mult_21_n264) );
  FA_X1 p9_mult_21_U108 ( .A(p9_mult_21_n275), .B(p9_mult_21_n385), .CI(
        p9_mult_21_n273), .CO(p9_mult_21_n261), .S(p9_mult_21_n262) );
  FA_X1 p9_mult_21_U107 ( .A(p9_mult_21_n264), .B(p9_mult_21_n266), .CI(
        p9_mult_21_n271), .CO(p9_mult_21_n259), .S(p9_mult_21_n260) );
  FA_X1 p9_mult_21_U106 ( .A(p9_mult_21_n262), .B(p9_mult_21_n269), .CI(
        p9_mult_21_n260), .CO(p9_mult_21_n257), .S(p9_mult_21_n258) );
  HA_X1 p9_mult_21_U105 ( .A(p9_mult_21_n317), .B(p9_mult_21_n336), .CO(
        p9_mult_21_n255), .S(p9_mult_21_n256) );
  FA_X1 p9_mult_21_U104 ( .A(p9_mult_21_n409), .B(p9_mult_21_n372), .CI(
        p9_mult_21_n396), .CO(p9_mult_21_n253), .S(p9_mult_21_n254) );
  FA_X1 p9_mult_21_U103 ( .A(p9_mult_21_n348), .B(p9_mult_21_n384), .CI(
        p9_mult_21_n360), .CO(p9_mult_21_n251), .S(p9_mult_21_n252) );
  FA_X1 p9_mult_21_U102 ( .A(p9_mult_21_n265), .B(p9_mult_21_n256), .CI(
        p9_mult_21_n263), .CO(p9_mult_21_n249), .S(p9_mult_21_n250) );
  FA_X1 p9_mult_21_U101 ( .A(p9_mult_21_n254), .B(p9_mult_21_n252), .CI(
        p9_mult_21_n261), .CO(p9_mult_21_n247), .S(p9_mult_21_n248) );
  FA_X1 p9_mult_21_U100 ( .A(p9_mult_21_n259), .B(p9_mult_21_n250), .CI(
        p9_mult_21_n248), .CO(p9_mult_21_n245), .S(p9_mult_21_n246) );
  FA_X1 p9_mult_21_U97 ( .A(p9_mult_21_n395), .B(p9_mult_21_n359), .CI(
        p9_mult_21_n408), .CO(p9_mult_21_n241), .S(p9_mult_21_n242) );
  FA_X1 p9_mult_21_U96 ( .A(p9_mult_21_n335), .B(p9_mult_21_n371), .CI(
        p9_mult_21_n255), .CO(p9_mult_21_n239), .S(p9_mult_21_n240) );
  FA_X1 p9_mult_21_U95 ( .A(p9_mult_21_n253), .B(p9_mult_21_n244), .CI(
        p9_mult_21_n251), .CO(p9_mult_21_n237), .S(p9_mult_21_n238) );
  FA_X1 p9_mult_21_U94 ( .A(p9_mult_21_n240), .B(p9_mult_21_n242), .CI(
        p9_mult_21_n249), .CO(p9_mult_21_n235), .S(p9_mult_21_n236) );
  FA_X1 p9_mult_21_U93 ( .A(p9_mult_21_n247), .B(p9_mult_21_n238), .CI(
        p9_mult_21_n236), .CO(p9_mult_21_n233), .S(p9_mult_21_n234) );
  FA_X1 p9_mult_21_U91 ( .A(p9_mult_21_n382), .B(p9_mult_21_n346), .CI(
        p9_mult_21_n232), .CO(p9_mult_21_n229), .S(p9_mult_21_n230) );
  FA_X1 p9_mult_21_U90 ( .A(p9_mult_21_n334), .B(p9_mult_21_n370), .CI(
        p9_mult_21_n358), .CO(p9_mult_21_n227), .S(p9_mult_21_n228) );
  FA_X1 p9_mult_21_U89 ( .A(p9_mult_21_n241), .B(p9_mult_21_n243), .CI(
        p9_mult_21_n239), .CO(p9_mult_21_n225), .S(p9_mult_21_n226) );
  FA_X1 p9_mult_21_U88 ( .A(p9_mult_21_n230), .B(p9_mult_21_n228), .CI(
        p9_mult_21_n237), .CO(p9_mult_21_n223), .S(p9_mult_21_n224) );
  FA_X1 p9_mult_21_U87 ( .A(p9_mult_21_n235), .B(p9_mult_21_n226), .CI(
        p9_mult_21_n224), .CO(p9_mult_21_n221), .S(p9_mult_21_n222) );
  FA_X1 p9_mult_21_U86 ( .A(p9_mult_21_n231), .B(p9_mult_21_n333), .CI(
        p9_mult_21_n394), .CO(p9_mult_21_n219), .S(p9_mult_21_n220) );
  FA_X1 p9_mult_21_U85 ( .A(p9_mult_21_n345), .B(p9_mult_21_n381), .CI(
        p9_mult_21_n357), .CO(p9_mult_21_n217), .S(p9_mult_21_n218) );
  FA_X1 p9_mult_21_U84 ( .A(p9_mult_21_n229), .B(p9_mult_21_n369), .CI(
        p9_mult_21_n227), .CO(p9_mult_21_n215), .S(p9_mult_21_n216) );
  FA_X1 p9_mult_21_U83 ( .A(p9_mult_21_n220), .B(p9_mult_21_n218), .CI(
        p9_mult_21_n225), .CO(p9_mult_21_n213), .S(p9_mult_21_n214) );
  FA_X1 p9_mult_21_U82 ( .A(p9_mult_21_n223), .B(p9_mult_21_n216), .CI(
        p9_mult_21_n214), .CO(p9_mult_21_n211), .S(p9_mult_21_n212) );
  FA_X1 p9_mult_21_U80 ( .A(p9_mult_21_n368), .B(p9_mult_21_n344), .CI(
        p9_mult_21_n210), .CO(p9_mult_21_n207), .S(p9_mult_21_n208) );
  FA_X1 p9_mult_21_U79 ( .A(p9_mult_21_n332), .B(p9_mult_21_n356), .CI(
        p9_mult_21_n219), .CO(p9_mult_21_n205), .S(p9_mult_21_n206) );
  FA_X1 p9_mult_21_U78 ( .A(p9_mult_21_n208), .B(p9_mult_21_n217), .CI(
        p9_mult_21_n215), .CO(p9_mult_21_n203), .S(p9_mult_21_n204) );
  FA_X1 p9_mult_21_U77 ( .A(p9_mult_21_n213), .B(p9_mult_21_n206), .CI(
        p9_mult_21_n204), .CO(p9_mult_21_n201), .S(p9_mult_21_n202) );
  FA_X1 p9_mult_21_U76 ( .A(p9_mult_21_n209), .B(p9_mult_21_n331), .CI(
        p9_mult_21_n380), .CO(p9_mult_21_n199), .S(p9_mult_21_n200) );
  FA_X1 p9_mult_21_U75 ( .A(p9_mult_21_n355), .B(p9_mult_21_n343), .CI(
        p9_mult_21_n367), .CO(p9_mult_21_n197), .S(p9_mult_21_n198) );
  FA_X1 p9_mult_21_U74 ( .A(p9_mult_21_n198), .B(p9_mult_21_n207), .CI(
        p9_mult_21_n200), .CO(p9_mult_21_n195), .S(p9_mult_21_n196) );
  FA_X1 p9_mult_21_U73 ( .A(p9_mult_21_n203), .B(p9_mult_21_n205), .CI(
        p9_mult_21_n196), .CO(p9_mult_21_n193), .S(p9_mult_21_n194) );
  FA_X1 p9_mult_21_U71 ( .A(p9_mult_21_n330), .B(p9_mult_21_n342), .CI(
        p9_mult_21_n192), .CO(p9_mult_21_n189), .S(p9_mult_21_n190) );
  FA_X1 p9_mult_21_U70 ( .A(p9_mult_21_n199), .B(p9_mult_21_n354), .CI(
        p9_mult_21_n197), .CO(p9_mult_21_n187), .S(p9_mult_21_n188) );
  FA_X1 p9_mult_21_U69 ( .A(p9_mult_21_n188), .B(p9_mult_21_n190), .CI(
        p9_mult_21_n195), .CO(p9_mult_21_n185), .S(p9_mult_21_n186) );
  FA_X1 p9_mult_21_U68 ( .A(p9_mult_21_n191), .B(p9_mult_21_n329), .CI(
        p9_mult_21_n366), .CO(p9_mult_21_n183), .S(p9_mult_21_n184) );
  FA_X1 p9_mult_21_U67 ( .A(p9_mult_21_n341), .B(p9_mult_21_n353), .CI(
        p9_mult_21_n189), .CO(p9_mult_21_n181), .S(p9_mult_21_n182) );
  FA_X1 p9_mult_21_U66 ( .A(p9_mult_21_n187), .B(p9_mult_21_n184), .CI(
        p9_mult_21_n182), .CO(p9_mult_21_n179), .S(p9_mult_21_n180) );
  FA_X1 p9_mult_21_U64 ( .A(p9_mult_21_n328), .B(p9_mult_21_n340), .CI(
        p9_mult_21_n178), .CO(p9_mult_21_n175), .S(p9_mult_21_n176) );
  FA_X1 p9_mult_21_U63 ( .A(p9_mult_21_n176), .B(p9_mult_21_n183), .CI(
        p9_mult_21_n181), .CO(p9_mult_21_n173), .S(p9_mult_21_n174) );
  FA_X1 p9_mult_21_U62 ( .A(p9_mult_21_n327), .B(p9_mult_21_n177), .CI(
        p9_mult_21_n352), .CO(p9_mult_21_n171), .S(p9_mult_21_n172) );
  FA_X1 p9_mult_21_U61 ( .A(p9_mult_21_n175), .B(p9_mult_21_n339), .CI(
        p9_mult_21_n172), .CO(p9_mult_21_n169), .S(p9_mult_21_n170) );
  FA_X1 p9_mult_21_U59 ( .A(p9_mult_21_n168), .B(p9_mult_21_n326), .CI(
        p9_mult_21_n171), .CO(p9_mult_21_n165), .S(p9_mult_21_n166) );
  FA_X1 p9_mult_21_U58 ( .A(p9_mult_21_n325), .B(p9_mult_21_n167), .CI(
        p9_mult_21_n338), .CO(p9_mult_21_n163), .S(p9_mult_21_n164) );
  FA_X1 p9_mult_21_U44 ( .A(p9_mult_21_n246), .B(p9_mult_21_n257), .CI(
        p9_mult_21_n149), .CO(p9_mult_21_n148), .S(temp4[0]) );
  FA_X1 p9_mult_21_U43 ( .A(p9_mult_21_n234), .B(p9_mult_21_n245), .CI(
        p9_mult_21_n148), .CO(p9_mult_21_n147), .S(temp4[1]) );
  FA_X1 p9_mult_21_U42 ( .A(p9_mult_21_n222), .B(p9_mult_21_n233), .CI(
        p9_mult_21_n147), .CO(p9_mult_21_n146), .S(temp4[2]) );
  FA_X1 p9_mult_21_U41 ( .A(p9_mult_21_n212), .B(p9_mult_21_n221), .CI(
        p9_mult_21_n146), .CO(p9_mult_21_n145), .S(temp4[3]) );
  FA_X1 p9_mult_21_U40 ( .A(p9_mult_21_n202), .B(p9_mult_21_n211), .CI(
        p9_mult_21_n145), .CO(p9_mult_21_n144), .S(temp4[4]) );
  FA_X1 p9_mult_21_U39 ( .A(p9_mult_21_n194), .B(p9_mult_21_n201), .CI(
        p9_mult_21_n144), .CO(p9_mult_21_n143), .S(temp4[5]) );
  FA_X1 p9_mult_21_U38 ( .A(p9_mult_21_n186), .B(p9_mult_21_n193), .CI(
        p9_mult_21_n143), .CO(p9_mult_21_n142), .S(temp4[6]) );
  FA_X1 p9_mult_21_U37 ( .A(p9_mult_21_n180), .B(p9_mult_21_n185), .CI(
        p9_mult_21_n142), .CO(p9_mult_21_n141), .S(temp4[7]) );
  FA_X1 p9_mult_21_U30 ( .A(p9_mult_21_n174), .B(p9_mult_21_n179), .CI(
        p9_mult_21_n141), .CO(p9_mult_21_n140), .S(temp4[8]) );
  FA_X1 p9_mult_21_U20 ( .A(p9_mult_21_n170), .B(p9_mult_21_n173), .CI(
        p9_mult_21_n140), .CO(p9_mult_21_n139), .S(temp4[9]) );
  FA_X1 p9_mult_21_U10 ( .A(p9_mult_21_n166), .B(p9_mult_21_n169), .CI(
        p9_mult_21_n139), .CO(p9_mult_21_n138), .S(temp4[10]) );
  FA_X1 p9_mult_21_U9 ( .A(p9_mult_21_n165), .B(p9_mult_21_n164), .CI(
        p9_mult_21_n138), .CO(p9_mult_21_n137), .S(temp4[11]) );
  FA_X1 p9_mult_21_U8 ( .A(p9_mult_21_n163), .B(p9_mult_21_n162), .CI(
        p9_mult_21_n137), .CO(p9_mult_21_n136), .S(temp4[12]) );
  NAND2_X1 REG4_1_U34 ( .A1(temp4[4]), .A2(REG4_1_n43), .ZN(REG4_1_n85) );
  OAI21_X1 REG4_1_U33 ( .B1(REG4_1_n45), .B2(REG4_1_n66), .A(REG4_1_n85), .ZN(
        REG4_1_n57) );
  NAND2_X1 REG4_1_U32 ( .A1(temp4[3]), .A2(REG4_1_n43), .ZN(REG4_1_n86) );
  OAI21_X1 REG4_1_U31 ( .B1(REG4_1_n45), .B2(REG4_1_n65), .A(REG4_1_n86), .ZN(
        REG4_1_n58) );
  NAND2_X1 REG4_1_U30 ( .A1(temp4[2]), .A2(REG4_1_n43), .ZN(REG4_1_n87) );
  OAI21_X1 REG4_1_U29 ( .B1(REG4_1_n45), .B2(REG4_1_n64), .A(REG4_1_n87), .ZN(
        REG4_1_n59) );
  NAND2_X1 REG4_1_U28 ( .A1(temp4[5]), .A2(REG4_1_n43), .ZN(REG4_1_n84) );
  OAI21_X1 REG4_1_U27 ( .B1(REG4_1_n44), .B2(REG4_1_n67), .A(REG4_1_n84), .ZN(
        REG4_1_n56) );
  NAND2_X1 REG4_1_U26 ( .A1(temp4[9]), .A2(REG4_1_n43), .ZN(REG4_1_n80) );
  OAI21_X1 REG4_1_U25 ( .B1(REG4_1_n44), .B2(REG4_1_n71), .A(REG4_1_n80), .ZN(
        REG4_1_n52) );
  NAND2_X1 REG4_1_U24 ( .A1(temp4[8]), .A2(REG4_1_n44), .ZN(REG4_1_n81) );
  OAI21_X1 REG4_1_U23 ( .B1(REG4_1_n44), .B2(REG4_1_n70), .A(REG4_1_n81), .ZN(
        REG4_1_n53) );
  NAND2_X1 REG4_1_U22 ( .A1(temp4[7]), .A2(REG4_1_n43), .ZN(REG4_1_n82) );
  OAI21_X1 REG4_1_U21 ( .B1(REG4_1_n44), .B2(REG4_1_n69), .A(REG4_1_n82), .ZN(
        REG4_1_n54) );
  NAND2_X1 REG4_1_U20 ( .A1(temp4[6]), .A2(REG4_1_n43), .ZN(REG4_1_n83) );
  OAI21_X1 REG4_1_U19 ( .B1(REG4_1_n44), .B2(REG4_1_n68), .A(REG4_1_n83), .ZN(
        REG4_1_n55) );
  NAND2_X1 REG4_1_U18 ( .A1(temp4[1]), .A2(REG4_1_n43), .ZN(REG4_1_n88) );
  OAI21_X1 REG4_1_U17 ( .B1(REG4_1_n44), .B2(REG4_1_n63), .A(REG4_1_n88), .ZN(
        REG4_1_n60) );
  NAND2_X1 REG4_1_U16 ( .A1(temp4[0]), .A2(REG4_1_n43), .ZN(REG4_1_n89) );
  OAI21_X1 REG4_1_U15 ( .B1(REG4_1_n44), .B2(REG4_1_n62), .A(REG4_1_n89), .ZN(
        REG4_1_n61) );
  NAND2_X1 REG4_1_U14 ( .A1(temp4[10]), .A2(REG4_1_n44), .ZN(REG4_1_n79) );
  OAI21_X1 REG4_1_U13 ( .B1(REG4_1_n44), .B2(REG4_1_n72), .A(REG4_1_n79), .ZN(
        REG4_1_n51) );
  NAND2_X1 REG4_1_U12 ( .A1(temp4[12]), .A2(REG4_1_n43), .ZN(REG4_1_n77) );
  OAI21_X1 REG4_1_U11 ( .B1(REG4_1_n44), .B2(REG4_1_n74), .A(REG4_1_n77), .ZN(
        REG4_1_n49) );
  NAND2_X1 REG4_1_U10 ( .A1(temp4[11]), .A2(REG4_1_n43), .ZN(REG4_1_n78) );
  OAI21_X1 REG4_1_U9 ( .B1(REG4_1_n44), .B2(REG4_1_n73), .A(REG4_1_n78), .ZN(
        REG4_1_n50) );
  NAND2_X1 REG4_1_U8 ( .A1(temp4[13]), .A2(REG4_1_n43), .ZN(REG4_1_n76) );
  OAI21_X1 REG4_1_U7 ( .B1(REG4_1_n44), .B2(REG4_1_n75), .A(REG4_1_n76), .ZN(
        REG4_1_n48) );
  BUF_X1 REG4_1_U6 ( .A(n47), .Z(REG4_1_n47) );
  BUF_X1 REG4_1_U5 ( .A(n47), .Z(REG4_1_n46) );
  BUF_X1 REG4_1_U4 ( .A(VIN), .Z(REG4_1_n45) );
  BUF_X1 REG4_1_U3 ( .A(VIN), .Z(REG4_1_n43) );
  BUF_X1 REG4_1_U2 ( .A(VIN), .Z(REG4_1_n44) );
  DFFR_X1 REG4_1_q_reg_0_ ( .D(REG4_1_n61), .CK(CLK), .RN(REG4_1_n47), .Q(
        mul4_reg[0]), .QN(REG4_1_n62) );
  DFFR_X1 REG4_1_q_reg_1_ ( .D(REG4_1_n60), .CK(CLK), .RN(REG4_1_n47), .Q(
        mul4_reg[1]), .QN(REG4_1_n63) );
  DFFR_X1 REG4_1_q_reg_2_ ( .D(REG4_1_n59), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[2]), .QN(REG4_1_n64) );
  DFFR_X1 REG4_1_q_reg_3_ ( .D(REG4_1_n58), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[3]), .QN(REG4_1_n65) );
  DFFR_X1 REG4_1_q_reg_4_ ( .D(REG4_1_n57), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[4]), .QN(REG4_1_n66) );
  DFFR_X1 REG4_1_q_reg_5_ ( .D(REG4_1_n56), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[5]), .QN(REG4_1_n67) );
  DFFR_X1 REG4_1_q_reg_6_ ( .D(REG4_1_n55), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[6]), .QN(REG4_1_n68) );
  DFFR_X1 REG4_1_q_reg_7_ ( .D(REG4_1_n54), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[7]), .QN(REG4_1_n69) );
  DFFR_X1 REG4_1_q_reg_8_ ( .D(REG4_1_n53), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[8]), .QN(REG4_1_n70) );
  DFFR_X1 REG4_1_q_reg_9_ ( .D(REG4_1_n52), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[9]), .QN(REG4_1_n71) );
  DFFR_X1 REG4_1_q_reg_10_ ( .D(REG4_1_n51), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[10]), .QN(REG4_1_n72) );
  DFFR_X1 REG4_1_q_reg_11_ ( .D(REG4_1_n50), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[11]), .QN(REG4_1_n73) );
  DFFR_X1 REG4_1_q_reg_12_ ( .D(REG4_1_n49), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[12]), .QN(REG4_1_n74) );
  DFFR_X1 REG4_1_q_reg_13_ ( .D(REG4_1_n48), .CK(CLK), .RN(REG4_1_n46), .Q(
        mul4_reg[13]), .QN(REG4_1_n75) );
  XOR2_X1 p11_mult_21_U691 ( .A(reg2[2]), .B(reg2[1]), .Z(p11_mult_21_n798) );
  INV_X1 p11_mult_21_U690 ( .A(reg2[1]), .ZN(p11_mult_21_n655) );
  NOR2_X1 p11_mult_21_U689 ( .A1(p11_mult_21_n655), .A2(A1[1]), .ZN(
        p11_mult_21_n803) );
  INV_X1 p11_mult_21_U688 ( .A(p11_mult_21_n803), .ZN(p11_mult_21_n805) );
  NAND2_X1 p11_mult_21_U687 ( .A1(reg2[1]), .A2(p11_mult_21_n643), .ZN(
        p11_mult_21_n641) );
  XNOR2_X1 p11_mult_21_U686 ( .A(A1[2]), .B(reg2[1]), .ZN(p11_mult_21_n640) );
  OAI22_X1 p11_mult_21_U685 ( .A1(p11_mult_21_n805), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n640), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n804) );
  NAND2_X1 p11_mult_21_U684 ( .A1(p11_mult_21_n798), .A2(p11_mult_21_n804), 
        .ZN(p11_mult_21_n801) );
  NAND2_X1 p11_mult_21_U683 ( .A1(p11_mult_21_n803), .A2(p11_mult_21_n804), 
        .ZN(p11_mult_21_n802) );
  INV_X1 p11_mult_21_U682 ( .A(A1[0]), .ZN(p11_mult_21_n673) );
  MUX2_X1 p11_mult_21_U681 ( .A(p11_mult_21_n801), .B(p11_mult_21_n802), .S(
        p11_mult_21_n673), .Z(p11_mult_21_n800) );
  INV_X1 p11_mult_21_U680 ( .A(p11_mult_21_n800), .ZN(p11_mult_21_n795) );
  INV_X1 p11_mult_21_U679 ( .A(reg2[3]), .ZN(p11_mult_21_n771) );
  XNOR2_X1 p11_mult_21_U678 ( .A(p11_mult_21_n771), .B(reg2[2]), .ZN(
        p11_mult_21_n799) );
  NAND2_X1 p11_mult_21_U677 ( .A1(p11_mult_21_n658), .A2(p11_mult_21_n799), 
        .ZN(p11_mult_21_n657) );
  NAND3_X1 p11_mult_21_U676 ( .A1(p11_mult_21_n798), .A2(p11_mult_21_n673), 
        .A3(reg2[3]), .ZN(p11_mult_21_n797) );
  OAI21_X1 p11_mult_21_U675 ( .B1(p11_mult_21_n771), .B2(p11_mult_21_n657), 
        .A(p11_mult_21_n797), .ZN(p11_mult_21_n796) );
  AOI222_X1 p11_mult_21_U674 ( .A1(p11_mult_21_n795), .A2(p11_mult_21_n316), 
        .B1(p11_mult_21_n796), .B2(p11_mult_21_n795), .C1(p11_mult_21_n796), 
        .C2(p11_mult_21_n316), .ZN(p11_mult_21_n794) );
  INV_X1 p11_mult_21_U673 ( .A(p11_mult_21_n794), .ZN(p11_mult_21_n793) );
  AOI222_X1 p11_mult_21_U672 ( .A1(p11_mult_21_n793), .A2(p11_mult_21_n314), 
        .B1(p11_mult_21_n793), .B2(p11_mult_21_n315), .C1(p11_mult_21_n315), 
        .C2(p11_mult_21_n314), .ZN(p11_mult_21_n792) );
  INV_X1 p11_mult_21_U671 ( .A(p11_mult_21_n792), .ZN(p11_mult_21_n791) );
  AOI222_X1 p11_mult_21_U670 ( .A1(p11_mult_21_n791), .A2(p11_mult_21_n310), 
        .B1(p11_mult_21_n791), .B2(p11_mult_21_n313), .C1(p11_mult_21_n313), 
        .C2(p11_mult_21_n310), .ZN(p11_mult_21_n790) );
  INV_X1 p11_mult_21_U669 ( .A(p11_mult_21_n790), .ZN(p11_mult_21_n789) );
  AOI222_X1 p11_mult_21_U668 ( .A1(p11_mult_21_n789), .A2(p11_mult_21_n306), 
        .B1(p11_mult_21_n789), .B2(p11_mult_21_n309), .C1(p11_mult_21_n309), 
        .C2(p11_mult_21_n306), .ZN(p11_mult_21_n788) );
  INV_X1 p11_mult_21_U667 ( .A(p11_mult_21_n788), .ZN(p11_mult_21_n787) );
  AOI222_X1 p11_mult_21_U666 ( .A1(p11_mult_21_n787), .A2(p11_mult_21_n300), 
        .B1(p11_mult_21_n787), .B2(p11_mult_21_n305), .C1(p11_mult_21_n305), 
        .C2(p11_mult_21_n300), .ZN(p11_mult_21_n786) );
  INV_X1 p11_mult_21_U665 ( .A(p11_mult_21_n786), .ZN(p11_mult_21_n785) );
  AOI222_X1 p11_mult_21_U664 ( .A1(p11_mult_21_n785), .A2(p11_mult_21_n294), 
        .B1(p11_mult_21_n785), .B2(p11_mult_21_n299), .C1(p11_mult_21_n299), 
        .C2(p11_mult_21_n294), .ZN(p11_mult_21_n784) );
  INV_X1 p11_mult_21_U663 ( .A(p11_mult_21_n784), .ZN(p11_mult_21_n783) );
  AOI222_X1 p11_mult_21_U662 ( .A1(p11_mult_21_n783), .A2(p11_mult_21_n286), 
        .B1(p11_mult_21_n783), .B2(p11_mult_21_n293), .C1(p11_mult_21_n293), 
        .C2(p11_mult_21_n286), .ZN(p11_mult_21_n780) );
  INV_X1 p11_mult_21_U661 ( .A(p11_mult_21_n278), .ZN(p11_mult_21_n781) );
  INV_X1 p11_mult_21_U660 ( .A(p11_mult_21_n285), .ZN(p11_mult_21_n782) );
  OAI222_X1 p11_mult_21_U659 ( .A1(p11_mult_21_n780), .A2(p11_mult_21_n781), 
        .B1(p11_mult_21_n780), .B2(p11_mult_21_n782), .C1(p11_mult_21_n782), 
        .C2(p11_mult_21_n781), .ZN(p11_mult_21_n779) );
  AOI222_X1 p11_mult_21_U658 ( .A1(p11_mult_21_n779), .A2(p11_mult_21_n268), 
        .B1(p11_mult_21_n779), .B2(p11_mult_21_n277), .C1(p11_mult_21_n277), 
        .C2(p11_mult_21_n268), .ZN(p11_mult_21_n776) );
  INV_X1 p11_mult_21_U657 ( .A(p11_mult_21_n258), .ZN(p11_mult_21_n777) );
  INV_X1 p11_mult_21_U656 ( .A(p11_mult_21_n267), .ZN(p11_mult_21_n778) );
  OAI222_X1 p11_mult_21_U655 ( .A1(p11_mult_21_n776), .A2(p11_mult_21_n777), 
        .B1(p11_mult_21_n776), .B2(p11_mult_21_n778), .C1(p11_mult_21_n778), 
        .C2(p11_mult_21_n777), .ZN(p11_mult_21_n149) );
  XOR2_X1 p11_mult_21_U654 ( .A(A1[12]), .B(reg2[13]), .Z(p11_mult_21_n757) );
  INV_X1 p11_mult_21_U653 ( .A(reg2[11]), .ZN(p11_mult_21_n764) );
  INV_X1 p11_mult_21_U652 ( .A(reg2[13]), .ZN(p11_mult_21_n766) );
  XNOR2_X1 p11_mult_21_U651 ( .A(p11_mult_21_n766), .B(reg2[12]), .ZN(
        p11_mult_21_n775) );
  NAND2_X1 p11_mult_21_U650 ( .A1(p11_mult_21_n742), .A2(p11_mult_21_n775), 
        .ZN(p11_mult_21_n744) );
  INV_X1 p11_mult_21_U649 ( .A(p11_mult_21_n744), .ZN(p11_mult_21_n637) );
  INV_X1 p11_mult_21_U648 ( .A(p11_mult_21_n742), .ZN(p11_mult_21_n638) );
  XNOR2_X1 p11_mult_21_U647 ( .A(A1[13]), .B(p11_mult_21_n766), .ZN(
        p11_mult_21_n639) );
  AOI22_X1 p11_mult_21_U646 ( .A1(p11_mult_21_n757), .A2(p11_mult_21_n637), 
        .B1(p11_mult_21_n638), .B2(p11_mult_21_n639), .ZN(p11_mult_21_n162) );
  XNOR2_X1 p11_mult_21_U645 ( .A(A1[12]), .B(reg2[11]), .ZN(p11_mult_21_n739)
         );
  INV_X1 p11_mult_21_U644 ( .A(reg2[9]), .ZN(p11_mult_21_n762) );
  XNOR2_X1 p11_mult_21_U643 ( .A(p11_mult_21_n764), .B(reg2[10]), .ZN(
        p11_mult_21_n774) );
  NAND2_X1 p11_mult_21_U642 ( .A1(p11_mult_21_n725), .A2(p11_mult_21_n774), 
        .ZN(p11_mult_21_n727) );
  XNOR2_X1 p11_mult_21_U641 ( .A(A1[13]), .B(reg2[11]), .ZN(p11_mult_21_n741)
         );
  OAI22_X1 p11_mult_21_U640 ( .A1(p11_mult_21_n739), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n741), .ZN(p11_mult_21_n167) );
  INV_X1 p11_mult_21_U639 ( .A(p11_mult_21_n167), .ZN(p11_mult_21_n168) );
  XNOR2_X1 p11_mult_21_U638 ( .A(A1[12]), .B(reg2[9]), .ZN(p11_mult_21_n722)
         );
  INV_X1 p11_mult_21_U637 ( .A(reg2[7]), .ZN(p11_mult_21_n760) );
  XNOR2_X1 p11_mult_21_U636 ( .A(p11_mult_21_n762), .B(reg2[8]), .ZN(
        p11_mult_21_n773) );
  NAND2_X1 p11_mult_21_U635 ( .A1(p11_mult_21_n708), .A2(p11_mult_21_n773), 
        .ZN(p11_mult_21_n710) );
  XNOR2_X1 p11_mult_21_U634 ( .A(A1[13]), .B(reg2[9]), .ZN(p11_mult_21_n724)
         );
  OAI22_X1 p11_mult_21_U633 ( .A1(p11_mult_21_n722), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n724), .ZN(p11_mult_21_n177) );
  INV_X1 p11_mult_21_U632 ( .A(p11_mult_21_n177), .ZN(p11_mult_21_n178) );
  XNOR2_X1 p11_mult_21_U631 ( .A(A1[12]), .B(reg2[7]), .ZN(p11_mult_21_n705)
         );
  INV_X1 p11_mult_21_U630 ( .A(reg2[5]), .ZN(p11_mult_21_n758) );
  XNOR2_X1 p11_mult_21_U629 ( .A(p11_mult_21_n760), .B(reg2[6]), .ZN(
        p11_mult_21_n772) );
  NAND2_X1 p11_mult_21_U628 ( .A1(p11_mult_21_n691), .A2(p11_mult_21_n772), 
        .ZN(p11_mult_21_n693) );
  XNOR2_X1 p11_mult_21_U627 ( .A(A1[13]), .B(reg2[7]), .ZN(p11_mult_21_n707)
         );
  OAI22_X1 p11_mult_21_U626 ( .A1(p11_mult_21_n705), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n707), .ZN(p11_mult_21_n191) );
  INV_X1 p11_mult_21_U625 ( .A(p11_mult_21_n191), .ZN(p11_mult_21_n192) );
  XNOR2_X1 p11_mult_21_U624 ( .A(A1[12]), .B(reg2[5]), .ZN(p11_mult_21_n688)
         );
  XNOR2_X1 p11_mult_21_U623 ( .A(p11_mult_21_n758), .B(reg2[4]), .ZN(
        p11_mult_21_n770) );
  NAND2_X1 p11_mult_21_U622 ( .A1(p11_mult_21_n674), .A2(p11_mult_21_n770), 
        .ZN(p11_mult_21_n676) );
  XNOR2_X1 p11_mult_21_U621 ( .A(A1[13]), .B(reg2[5]), .ZN(p11_mult_21_n690)
         );
  OAI22_X1 p11_mult_21_U620 ( .A1(p11_mult_21_n688), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n690), .ZN(p11_mult_21_n209) );
  INV_X1 p11_mult_21_U619 ( .A(p11_mult_21_n209), .ZN(p11_mult_21_n210) );
  XNOR2_X1 p11_mult_21_U618 ( .A(A1[12]), .B(reg2[3]), .ZN(p11_mult_21_n670)
         );
  XNOR2_X1 p11_mult_21_U617 ( .A(A1[13]), .B(reg2[3]), .ZN(p11_mult_21_n672)
         );
  OAI22_X1 p11_mult_21_U616 ( .A1(p11_mult_21_n670), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n672), .ZN(p11_mult_21_n231) );
  INV_X1 p11_mult_21_U615 ( .A(p11_mult_21_n231), .ZN(p11_mult_21_n232) );
  XNOR2_X1 p11_mult_21_U614 ( .A(A1[3]), .B(reg2[11]), .ZN(p11_mult_21_n730)
         );
  XNOR2_X1 p11_mult_21_U613 ( .A(A1[4]), .B(reg2[11]), .ZN(p11_mult_21_n731)
         );
  OAI22_X1 p11_mult_21_U612 ( .A1(p11_mult_21_n730), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n731), .ZN(p11_mult_21_n768) );
  XNOR2_X1 p11_mult_21_U611 ( .A(A1[9]), .B(reg2[5]), .ZN(p11_mult_21_n685) );
  XNOR2_X1 p11_mult_21_U610 ( .A(A1[10]), .B(reg2[5]), .ZN(p11_mult_21_n686)
         );
  OAI22_X1 p11_mult_21_U609 ( .A1(p11_mult_21_n685), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n686), .ZN(p11_mult_21_n769) );
  OR2_X1 p11_mult_21_U608 ( .A1(p11_mult_21_n768), .A2(p11_mult_21_n769), .ZN(
        p11_mult_21_n243) );
  XNOR2_X1 p11_mult_21_U607 ( .A(p11_mult_21_n768), .B(p11_mult_21_n769), .ZN(
        p11_mult_21_n244) );
  NAND3_X1 p11_mult_21_U606 ( .A1(p11_mult_21_n638), .A2(p11_mult_21_n673), 
        .A3(reg2[13]), .ZN(p11_mult_21_n767) );
  OAI21_X1 p11_mult_21_U605 ( .B1(p11_mult_21_n766), .B2(p11_mult_21_n744), 
        .A(p11_mult_21_n767), .ZN(p11_mult_21_n317) );
  OR3_X1 p11_mult_21_U604 ( .A1(p11_mult_21_n725), .A2(A1[0]), .A3(
        p11_mult_21_n764), .ZN(p11_mult_21_n765) );
  OAI21_X1 p11_mult_21_U603 ( .B1(p11_mult_21_n764), .B2(p11_mult_21_n727), 
        .A(p11_mult_21_n765), .ZN(p11_mult_21_n318) );
  OR3_X1 p11_mult_21_U602 ( .A1(p11_mult_21_n708), .A2(A1[0]), .A3(
        p11_mult_21_n762), .ZN(p11_mult_21_n763) );
  OAI21_X1 p11_mult_21_U601 ( .B1(p11_mult_21_n762), .B2(p11_mult_21_n710), 
        .A(p11_mult_21_n763), .ZN(p11_mult_21_n319) );
  OR3_X1 p11_mult_21_U600 ( .A1(p11_mult_21_n691), .A2(A1[0]), .A3(
        p11_mult_21_n760), .ZN(p11_mult_21_n761) );
  OAI21_X1 p11_mult_21_U599 ( .B1(p11_mult_21_n760), .B2(p11_mult_21_n693), 
        .A(p11_mult_21_n761), .ZN(p11_mult_21_n320) );
  OR3_X1 p11_mult_21_U598 ( .A1(p11_mult_21_n674), .A2(A1[0]), .A3(
        p11_mult_21_n758), .ZN(p11_mult_21_n759) );
  OAI21_X1 p11_mult_21_U597 ( .B1(p11_mult_21_n758), .B2(p11_mult_21_n676), 
        .A(p11_mult_21_n759), .ZN(p11_mult_21_n321) );
  XNOR2_X1 p11_mult_21_U596 ( .A(A1[11]), .B(reg2[13]), .ZN(p11_mult_21_n755)
         );
  INV_X1 p11_mult_21_U595 ( .A(p11_mult_21_n757), .ZN(p11_mult_21_n756) );
  OAI22_X1 p11_mult_21_U594 ( .A1(p11_mult_21_n755), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n756), .ZN(p11_mult_21_n325) );
  XNOR2_X1 p11_mult_21_U593 ( .A(A1[10]), .B(reg2[13]), .ZN(p11_mult_21_n754)
         );
  OAI22_X1 p11_mult_21_U592 ( .A1(p11_mult_21_n754), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n755), .ZN(p11_mult_21_n326) );
  XNOR2_X1 p11_mult_21_U591 ( .A(A1[9]), .B(reg2[13]), .ZN(p11_mult_21_n753)
         );
  OAI22_X1 p11_mult_21_U590 ( .A1(p11_mult_21_n753), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n754), .ZN(p11_mult_21_n327) );
  XNOR2_X1 p11_mult_21_U589 ( .A(A1[8]), .B(reg2[13]), .ZN(p11_mult_21_n752)
         );
  OAI22_X1 p11_mult_21_U588 ( .A1(p11_mult_21_n752), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n753), .ZN(p11_mult_21_n328) );
  XNOR2_X1 p11_mult_21_U587 ( .A(A1[7]), .B(reg2[13]), .ZN(p11_mult_21_n751)
         );
  OAI22_X1 p11_mult_21_U586 ( .A1(p11_mult_21_n751), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n752), .ZN(p11_mult_21_n329) );
  XNOR2_X1 p11_mult_21_U585 ( .A(A1[6]), .B(reg2[13]), .ZN(p11_mult_21_n750)
         );
  OAI22_X1 p11_mult_21_U584 ( .A1(p11_mult_21_n750), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n751), .ZN(p11_mult_21_n330) );
  XNOR2_X1 p11_mult_21_U583 ( .A(A1[5]), .B(reg2[13]), .ZN(p11_mult_21_n749)
         );
  OAI22_X1 p11_mult_21_U582 ( .A1(p11_mult_21_n749), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n750), .ZN(p11_mult_21_n331) );
  XNOR2_X1 p11_mult_21_U581 ( .A(A1[4]), .B(reg2[13]), .ZN(p11_mult_21_n748)
         );
  OAI22_X1 p11_mult_21_U580 ( .A1(p11_mult_21_n748), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n749), .ZN(p11_mult_21_n332) );
  XNOR2_X1 p11_mult_21_U579 ( .A(A1[3]), .B(reg2[13]), .ZN(p11_mult_21_n747)
         );
  OAI22_X1 p11_mult_21_U578 ( .A1(p11_mult_21_n747), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n748), .ZN(p11_mult_21_n333) );
  XNOR2_X1 p11_mult_21_U577 ( .A(A1[2]), .B(reg2[13]), .ZN(p11_mult_21_n746)
         );
  OAI22_X1 p11_mult_21_U576 ( .A1(p11_mult_21_n746), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n747), .ZN(p11_mult_21_n334) );
  XNOR2_X1 p11_mult_21_U575 ( .A(A1[1]), .B(reg2[13]), .ZN(p11_mult_21_n745)
         );
  OAI22_X1 p11_mult_21_U574 ( .A1(p11_mult_21_n745), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n746), .ZN(p11_mult_21_n335) );
  XNOR2_X1 p11_mult_21_U573 ( .A(reg2[13]), .B(A1[0]), .ZN(p11_mult_21_n743)
         );
  OAI22_X1 p11_mult_21_U572 ( .A1(p11_mult_21_n743), .A2(p11_mult_21_n744), 
        .B1(p11_mult_21_n742), .B2(p11_mult_21_n745), .ZN(p11_mult_21_n336) );
  NOR2_X1 p11_mult_21_U571 ( .A1(p11_mult_21_n673), .A2(p11_mult_21_n742), 
        .ZN(p11_mult_21_n337) );
  AOI21_X1 p11_mult_21_U570 ( .B1(p11_mult_21_n727), .B2(p11_mult_21_n725), 
        .A(p11_mult_21_n741), .ZN(p11_mult_21_n740) );
  INV_X1 p11_mult_21_U569 ( .A(p11_mult_21_n740), .ZN(p11_mult_21_n338) );
  XNOR2_X1 p11_mult_21_U568 ( .A(A1[11]), .B(reg2[11]), .ZN(p11_mult_21_n738)
         );
  OAI22_X1 p11_mult_21_U567 ( .A1(p11_mult_21_n738), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n739), .ZN(p11_mult_21_n339) );
  XNOR2_X1 p11_mult_21_U566 ( .A(A1[10]), .B(reg2[11]), .ZN(p11_mult_21_n737)
         );
  OAI22_X1 p11_mult_21_U565 ( .A1(p11_mult_21_n737), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n738), .ZN(p11_mult_21_n340) );
  XNOR2_X1 p11_mult_21_U564 ( .A(A1[9]), .B(reg2[11]), .ZN(p11_mult_21_n736)
         );
  OAI22_X1 p11_mult_21_U563 ( .A1(p11_mult_21_n736), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n737), .ZN(p11_mult_21_n341) );
  XNOR2_X1 p11_mult_21_U562 ( .A(A1[8]), .B(reg2[11]), .ZN(p11_mult_21_n735)
         );
  OAI22_X1 p11_mult_21_U561 ( .A1(p11_mult_21_n735), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n736), .ZN(p11_mult_21_n342) );
  XNOR2_X1 p11_mult_21_U560 ( .A(A1[7]), .B(reg2[11]), .ZN(p11_mult_21_n734)
         );
  OAI22_X1 p11_mult_21_U559 ( .A1(p11_mult_21_n734), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n735), .ZN(p11_mult_21_n343) );
  XNOR2_X1 p11_mult_21_U558 ( .A(A1[6]), .B(reg2[11]), .ZN(p11_mult_21_n733)
         );
  OAI22_X1 p11_mult_21_U557 ( .A1(p11_mult_21_n733), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n734), .ZN(p11_mult_21_n344) );
  XNOR2_X1 p11_mult_21_U556 ( .A(A1[5]), .B(reg2[11]), .ZN(p11_mult_21_n732)
         );
  OAI22_X1 p11_mult_21_U555 ( .A1(p11_mult_21_n732), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n733), .ZN(p11_mult_21_n345) );
  OAI22_X1 p11_mult_21_U554 ( .A1(p11_mult_21_n731), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n732), .ZN(p11_mult_21_n346) );
  XNOR2_X1 p11_mult_21_U553 ( .A(A1[2]), .B(reg2[11]), .ZN(p11_mult_21_n729)
         );
  OAI22_X1 p11_mult_21_U552 ( .A1(p11_mult_21_n729), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n730), .ZN(p11_mult_21_n348) );
  XNOR2_X1 p11_mult_21_U551 ( .A(A1[1]), .B(reg2[11]), .ZN(p11_mult_21_n728)
         );
  OAI22_X1 p11_mult_21_U550 ( .A1(p11_mult_21_n728), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n729), .ZN(p11_mult_21_n349) );
  XNOR2_X1 p11_mult_21_U549 ( .A(reg2[11]), .B(A1[0]), .ZN(p11_mult_21_n726)
         );
  OAI22_X1 p11_mult_21_U548 ( .A1(p11_mult_21_n726), .A2(p11_mult_21_n727), 
        .B1(p11_mult_21_n725), .B2(p11_mult_21_n728), .ZN(p11_mult_21_n350) );
  NOR2_X1 p11_mult_21_U547 ( .A1(p11_mult_21_n673), .A2(p11_mult_21_n725), 
        .ZN(p11_mult_21_n351) );
  AOI21_X1 p11_mult_21_U546 ( .B1(p11_mult_21_n710), .B2(p11_mult_21_n708), 
        .A(p11_mult_21_n724), .ZN(p11_mult_21_n723) );
  INV_X1 p11_mult_21_U545 ( .A(p11_mult_21_n723), .ZN(p11_mult_21_n352) );
  XNOR2_X1 p11_mult_21_U544 ( .A(A1[11]), .B(reg2[9]), .ZN(p11_mult_21_n721)
         );
  OAI22_X1 p11_mult_21_U543 ( .A1(p11_mult_21_n721), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n722), .ZN(p11_mult_21_n353) );
  XNOR2_X1 p11_mult_21_U542 ( .A(A1[10]), .B(reg2[9]), .ZN(p11_mult_21_n720)
         );
  OAI22_X1 p11_mult_21_U541 ( .A1(p11_mult_21_n720), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n721), .ZN(p11_mult_21_n354) );
  XNOR2_X1 p11_mult_21_U540 ( .A(A1[9]), .B(reg2[9]), .ZN(p11_mult_21_n719) );
  OAI22_X1 p11_mult_21_U539 ( .A1(p11_mult_21_n719), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n720), .ZN(p11_mult_21_n355) );
  XNOR2_X1 p11_mult_21_U538 ( .A(A1[8]), .B(reg2[9]), .ZN(p11_mult_21_n718) );
  OAI22_X1 p11_mult_21_U537 ( .A1(p11_mult_21_n718), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n719), .ZN(p11_mult_21_n356) );
  XNOR2_X1 p11_mult_21_U536 ( .A(A1[7]), .B(reg2[9]), .ZN(p11_mult_21_n717) );
  OAI22_X1 p11_mult_21_U535 ( .A1(p11_mult_21_n717), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n718), .ZN(p11_mult_21_n357) );
  XNOR2_X1 p11_mult_21_U534 ( .A(A1[6]), .B(reg2[9]), .ZN(p11_mult_21_n716) );
  OAI22_X1 p11_mult_21_U533 ( .A1(p11_mult_21_n716), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n717), .ZN(p11_mult_21_n358) );
  XNOR2_X1 p11_mult_21_U532 ( .A(A1[5]), .B(reg2[9]), .ZN(p11_mult_21_n715) );
  OAI22_X1 p11_mult_21_U531 ( .A1(p11_mult_21_n715), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n716), .ZN(p11_mult_21_n359) );
  XNOR2_X1 p11_mult_21_U530 ( .A(A1[4]), .B(reg2[9]), .ZN(p11_mult_21_n714) );
  OAI22_X1 p11_mult_21_U529 ( .A1(p11_mult_21_n714), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n715), .ZN(p11_mult_21_n360) );
  XNOR2_X1 p11_mult_21_U528 ( .A(A1[3]), .B(reg2[9]), .ZN(p11_mult_21_n713) );
  OAI22_X1 p11_mult_21_U527 ( .A1(p11_mult_21_n713), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n714), .ZN(p11_mult_21_n361) );
  XNOR2_X1 p11_mult_21_U526 ( .A(A1[2]), .B(reg2[9]), .ZN(p11_mult_21_n712) );
  OAI22_X1 p11_mult_21_U525 ( .A1(p11_mult_21_n712), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n713), .ZN(p11_mult_21_n362) );
  XNOR2_X1 p11_mult_21_U524 ( .A(A1[1]), .B(reg2[9]), .ZN(p11_mult_21_n711) );
  OAI22_X1 p11_mult_21_U523 ( .A1(p11_mult_21_n711), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n712), .ZN(p11_mult_21_n363) );
  XNOR2_X1 p11_mult_21_U522 ( .A(reg2[9]), .B(A1[0]), .ZN(p11_mult_21_n709) );
  OAI22_X1 p11_mult_21_U521 ( .A1(p11_mult_21_n709), .A2(p11_mult_21_n710), 
        .B1(p11_mult_21_n708), .B2(p11_mult_21_n711), .ZN(p11_mult_21_n364) );
  NOR2_X1 p11_mult_21_U520 ( .A1(p11_mult_21_n673), .A2(p11_mult_21_n708), 
        .ZN(p11_mult_21_n365) );
  AOI21_X1 p11_mult_21_U519 ( .B1(p11_mult_21_n693), .B2(p11_mult_21_n691), 
        .A(p11_mult_21_n707), .ZN(p11_mult_21_n706) );
  INV_X1 p11_mult_21_U518 ( .A(p11_mult_21_n706), .ZN(p11_mult_21_n366) );
  XNOR2_X1 p11_mult_21_U517 ( .A(A1[11]), .B(reg2[7]), .ZN(p11_mult_21_n704)
         );
  OAI22_X1 p11_mult_21_U516 ( .A1(p11_mult_21_n704), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n705), .ZN(p11_mult_21_n367) );
  XNOR2_X1 p11_mult_21_U515 ( .A(A1[10]), .B(reg2[7]), .ZN(p11_mult_21_n703)
         );
  OAI22_X1 p11_mult_21_U514 ( .A1(p11_mult_21_n703), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n704), .ZN(p11_mult_21_n368) );
  XNOR2_X1 p11_mult_21_U513 ( .A(A1[9]), .B(reg2[7]), .ZN(p11_mult_21_n702) );
  OAI22_X1 p11_mult_21_U512 ( .A1(p11_mult_21_n702), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n703), .ZN(p11_mult_21_n369) );
  XNOR2_X1 p11_mult_21_U511 ( .A(A1[8]), .B(reg2[7]), .ZN(p11_mult_21_n701) );
  OAI22_X1 p11_mult_21_U510 ( .A1(p11_mult_21_n701), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n702), .ZN(p11_mult_21_n370) );
  XNOR2_X1 p11_mult_21_U509 ( .A(A1[7]), .B(reg2[7]), .ZN(p11_mult_21_n700) );
  OAI22_X1 p11_mult_21_U508 ( .A1(p11_mult_21_n700), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n701), .ZN(p11_mult_21_n371) );
  XNOR2_X1 p11_mult_21_U507 ( .A(A1[6]), .B(reg2[7]), .ZN(p11_mult_21_n699) );
  OAI22_X1 p11_mult_21_U506 ( .A1(p11_mult_21_n699), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n700), .ZN(p11_mult_21_n372) );
  XNOR2_X1 p11_mult_21_U505 ( .A(A1[5]), .B(reg2[7]), .ZN(p11_mult_21_n698) );
  OAI22_X1 p11_mult_21_U504 ( .A1(p11_mult_21_n698), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n699), .ZN(p11_mult_21_n373) );
  XNOR2_X1 p11_mult_21_U503 ( .A(A1[4]), .B(reg2[7]), .ZN(p11_mult_21_n697) );
  OAI22_X1 p11_mult_21_U502 ( .A1(p11_mult_21_n697), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n698), .ZN(p11_mult_21_n374) );
  XNOR2_X1 p11_mult_21_U501 ( .A(A1[3]), .B(reg2[7]), .ZN(p11_mult_21_n696) );
  OAI22_X1 p11_mult_21_U500 ( .A1(p11_mult_21_n696), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n697), .ZN(p11_mult_21_n375) );
  XNOR2_X1 p11_mult_21_U499 ( .A(A1[2]), .B(reg2[7]), .ZN(p11_mult_21_n695) );
  OAI22_X1 p11_mult_21_U498 ( .A1(p11_mult_21_n695), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n696), .ZN(p11_mult_21_n376) );
  XNOR2_X1 p11_mult_21_U497 ( .A(A1[1]), .B(reg2[7]), .ZN(p11_mult_21_n694) );
  OAI22_X1 p11_mult_21_U496 ( .A1(p11_mult_21_n694), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n695), .ZN(p11_mult_21_n377) );
  XNOR2_X1 p11_mult_21_U495 ( .A(reg2[7]), .B(A1[0]), .ZN(p11_mult_21_n692) );
  OAI22_X1 p11_mult_21_U494 ( .A1(p11_mult_21_n692), .A2(p11_mult_21_n693), 
        .B1(p11_mult_21_n691), .B2(p11_mult_21_n694), .ZN(p11_mult_21_n378) );
  NOR2_X1 p11_mult_21_U493 ( .A1(p11_mult_21_n673), .A2(p11_mult_21_n691), 
        .ZN(p11_mult_21_n379) );
  AOI21_X1 p11_mult_21_U492 ( .B1(p11_mult_21_n676), .B2(p11_mult_21_n674), 
        .A(p11_mult_21_n690), .ZN(p11_mult_21_n689) );
  INV_X1 p11_mult_21_U491 ( .A(p11_mult_21_n689), .ZN(p11_mult_21_n380) );
  XNOR2_X1 p11_mult_21_U490 ( .A(A1[11]), .B(reg2[5]), .ZN(p11_mult_21_n687)
         );
  OAI22_X1 p11_mult_21_U489 ( .A1(p11_mult_21_n687), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n688), .ZN(p11_mult_21_n381) );
  OAI22_X1 p11_mult_21_U488 ( .A1(p11_mult_21_n686), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n687), .ZN(p11_mult_21_n382) );
  XNOR2_X1 p11_mult_21_U487 ( .A(A1[8]), .B(reg2[5]), .ZN(p11_mult_21_n684) );
  OAI22_X1 p11_mult_21_U486 ( .A1(p11_mult_21_n684), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n685), .ZN(p11_mult_21_n384) );
  XNOR2_X1 p11_mult_21_U485 ( .A(A1[7]), .B(reg2[5]), .ZN(p11_mult_21_n683) );
  OAI22_X1 p11_mult_21_U484 ( .A1(p11_mult_21_n683), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n684), .ZN(p11_mult_21_n385) );
  XNOR2_X1 p11_mult_21_U483 ( .A(A1[6]), .B(reg2[5]), .ZN(p11_mult_21_n682) );
  OAI22_X1 p11_mult_21_U482 ( .A1(p11_mult_21_n682), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n683), .ZN(p11_mult_21_n386) );
  XNOR2_X1 p11_mult_21_U481 ( .A(A1[5]), .B(reg2[5]), .ZN(p11_mult_21_n681) );
  OAI22_X1 p11_mult_21_U480 ( .A1(p11_mult_21_n681), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n682), .ZN(p11_mult_21_n387) );
  XNOR2_X1 p11_mult_21_U479 ( .A(A1[4]), .B(reg2[5]), .ZN(p11_mult_21_n680) );
  OAI22_X1 p11_mult_21_U478 ( .A1(p11_mult_21_n680), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n681), .ZN(p11_mult_21_n388) );
  XNOR2_X1 p11_mult_21_U477 ( .A(A1[3]), .B(reg2[5]), .ZN(p11_mult_21_n679) );
  OAI22_X1 p11_mult_21_U476 ( .A1(p11_mult_21_n679), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n680), .ZN(p11_mult_21_n389) );
  XNOR2_X1 p11_mult_21_U475 ( .A(A1[2]), .B(reg2[5]), .ZN(p11_mult_21_n678) );
  OAI22_X1 p11_mult_21_U474 ( .A1(p11_mult_21_n678), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n679), .ZN(p11_mult_21_n390) );
  XNOR2_X1 p11_mult_21_U473 ( .A(A1[1]), .B(reg2[5]), .ZN(p11_mult_21_n677) );
  OAI22_X1 p11_mult_21_U472 ( .A1(p11_mult_21_n677), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n678), .ZN(p11_mult_21_n391) );
  XNOR2_X1 p11_mult_21_U471 ( .A(reg2[5]), .B(A1[0]), .ZN(p11_mult_21_n675) );
  OAI22_X1 p11_mult_21_U470 ( .A1(p11_mult_21_n675), .A2(p11_mult_21_n676), 
        .B1(p11_mult_21_n674), .B2(p11_mult_21_n677), .ZN(p11_mult_21_n392) );
  NOR2_X1 p11_mult_21_U469 ( .A1(p11_mult_21_n673), .A2(p11_mult_21_n674), 
        .ZN(p11_mult_21_n393) );
  AOI21_X1 p11_mult_21_U468 ( .B1(p11_mult_21_n657), .B2(p11_mult_21_n658), 
        .A(p11_mult_21_n672), .ZN(p11_mult_21_n671) );
  INV_X1 p11_mult_21_U467 ( .A(p11_mult_21_n671), .ZN(p11_mult_21_n394) );
  XNOR2_X1 p11_mult_21_U466 ( .A(A1[11]), .B(reg2[3]), .ZN(p11_mult_21_n669)
         );
  OAI22_X1 p11_mult_21_U465 ( .A1(p11_mult_21_n669), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n670), .ZN(p11_mult_21_n395) );
  XNOR2_X1 p11_mult_21_U464 ( .A(A1[10]), .B(reg2[3]), .ZN(p11_mult_21_n668)
         );
  OAI22_X1 p11_mult_21_U463 ( .A1(p11_mult_21_n668), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n669), .ZN(p11_mult_21_n396) );
  XNOR2_X1 p11_mult_21_U462 ( .A(A1[9]), .B(reg2[3]), .ZN(p11_mult_21_n667) );
  OAI22_X1 p11_mult_21_U461 ( .A1(p11_mult_21_n667), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n668), .ZN(p11_mult_21_n397) );
  XNOR2_X1 p11_mult_21_U460 ( .A(A1[8]), .B(reg2[3]), .ZN(p11_mult_21_n666) );
  OAI22_X1 p11_mult_21_U459 ( .A1(p11_mult_21_n666), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n667), .ZN(p11_mult_21_n398) );
  XNOR2_X1 p11_mult_21_U458 ( .A(A1[7]), .B(reg2[3]), .ZN(p11_mult_21_n665) );
  OAI22_X1 p11_mult_21_U457 ( .A1(p11_mult_21_n665), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n666), .ZN(p11_mult_21_n399) );
  XNOR2_X1 p11_mult_21_U456 ( .A(A1[6]), .B(reg2[3]), .ZN(p11_mult_21_n664) );
  OAI22_X1 p11_mult_21_U455 ( .A1(p11_mult_21_n664), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n665), .ZN(p11_mult_21_n400) );
  XNOR2_X1 p11_mult_21_U454 ( .A(A1[5]), .B(reg2[3]), .ZN(p11_mult_21_n663) );
  OAI22_X1 p11_mult_21_U453 ( .A1(p11_mult_21_n663), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n664), .ZN(p11_mult_21_n401) );
  XNOR2_X1 p11_mult_21_U452 ( .A(A1[4]), .B(reg2[3]), .ZN(p11_mult_21_n662) );
  OAI22_X1 p11_mult_21_U451 ( .A1(p11_mult_21_n662), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n663), .ZN(p11_mult_21_n402) );
  XNOR2_X1 p11_mult_21_U450 ( .A(A1[3]), .B(reg2[3]), .ZN(p11_mult_21_n661) );
  OAI22_X1 p11_mult_21_U449 ( .A1(p11_mult_21_n661), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n662), .ZN(p11_mult_21_n403) );
  XNOR2_X1 p11_mult_21_U448 ( .A(A1[2]), .B(reg2[3]), .ZN(p11_mult_21_n660) );
  OAI22_X1 p11_mult_21_U447 ( .A1(p11_mult_21_n660), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n661), .ZN(p11_mult_21_n404) );
  XNOR2_X1 p11_mult_21_U446 ( .A(A1[1]), .B(reg2[3]), .ZN(p11_mult_21_n659) );
  OAI22_X1 p11_mult_21_U445 ( .A1(p11_mult_21_n659), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n660), .ZN(p11_mult_21_n405) );
  XNOR2_X1 p11_mult_21_U444 ( .A(reg2[3]), .B(A1[0]), .ZN(p11_mult_21_n656) );
  OAI22_X1 p11_mult_21_U443 ( .A1(p11_mult_21_n656), .A2(p11_mult_21_n657), 
        .B1(p11_mult_21_n658), .B2(p11_mult_21_n659), .ZN(p11_mult_21_n406) );
  XOR2_X1 p11_mult_21_U442 ( .A(A1[13]), .B(p11_mult_21_n655), .Z(
        p11_mult_21_n653) );
  AOI21_X1 p11_mult_21_U441 ( .B1(p11_mult_21_n641), .B2(p11_mult_21_n643), 
        .A(p11_mult_21_n653), .ZN(p11_mult_21_n654) );
  INV_X1 p11_mult_21_U440 ( .A(p11_mult_21_n654), .ZN(p11_mult_21_n408) );
  XNOR2_X1 p11_mult_21_U439 ( .A(A1[12]), .B(reg2[1]), .ZN(p11_mult_21_n652)
         );
  OAI22_X1 p11_mult_21_U438 ( .A1(p11_mult_21_n652), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n653), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n409) );
  XNOR2_X1 p11_mult_21_U437 ( .A(A1[11]), .B(reg2[1]), .ZN(p11_mult_21_n651)
         );
  OAI22_X1 p11_mult_21_U436 ( .A1(p11_mult_21_n651), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n652), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n410) );
  XNOR2_X1 p11_mult_21_U435 ( .A(A1[10]), .B(reg2[1]), .ZN(p11_mult_21_n650)
         );
  OAI22_X1 p11_mult_21_U434 ( .A1(p11_mult_21_n650), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n651), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n411) );
  XNOR2_X1 p11_mult_21_U433 ( .A(A1[9]), .B(reg2[1]), .ZN(p11_mult_21_n649) );
  OAI22_X1 p11_mult_21_U432 ( .A1(p11_mult_21_n649), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n650), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n412) );
  XNOR2_X1 p11_mult_21_U431 ( .A(A1[8]), .B(reg2[1]), .ZN(p11_mult_21_n648) );
  OAI22_X1 p11_mult_21_U430 ( .A1(p11_mult_21_n648), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n649), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n413) );
  XNOR2_X1 p11_mult_21_U429 ( .A(A1[7]), .B(reg2[1]), .ZN(p11_mult_21_n647) );
  OAI22_X1 p11_mult_21_U428 ( .A1(p11_mult_21_n647), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n648), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n414) );
  XNOR2_X1 p11_mult_21_U427 ( .A(A1[6]), .B(reg2[1]), .ZN(p11_mult_21_n646) );
  OAI22_X1 p11_mult_21_U426 ( .A1(p11_mult_21_n646), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n647), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n415) );
  XNOR2_X1 p11_mult_21_U425 ( .A(A1[5]), .B(reg2[1]), .ZN(p11_mult_21_n645) );
  OAI22_X1 p11_mult_21_U424 ( .A1(p11_mult_21_n645), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n646), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n416) );
  XNOR2_X1 p11_mult_21_U423 ( .A(A1[4]), .B(reg2[1]), .ZN(p11_mult_21_n644) );
  OAI22_X1 p11_mult_21_U422 ( .A1(p11_mult_21_n644), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n645), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n417) );
  XNOR2_X1 p11_mult_21_U421 ( .A(A1[3]), .B(reg2[1]), .ZN(p11_mult_21_n642) );
  OAI22_X1 p11_mult_21_U420 ( .A1(p11_mult_21_n642), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n644), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n418) );
  OAI22_X1 p11_mult_21_U419 ( .A1(p11_mult_21_n640), .A2(p11_mult_21_n641), 
        .B1(p11_mult_21_n642), .B2(p11_mult_21_n643), .ZN(p11_mult_21_n419) );
  OAI21_X1 p11_mult_21_U418 ( .B1(p11_mult_21_n637), .B2(p11_mult_21_n638), 
        .A(p11_mult_21_n639), .ZN(p11_mult_21_n636) );
  XOR2_X1 p11_mult_21_U417 ( .A(p11_mult_21_n636), .B(p11_mult_21_n136), .Z(
        p11_mult_21_n635) );
  XNOR2_X1 p11_mult_21_U416 ( .A(p11_mult_21_n162), .B(p11_mult_21_n635), .ZN(
        temp6[13]) );
  XOR2_X2 p11_mult_21_U415 ( .A(reg2[12]), .B(p11_mult_21_n764), .Z(
        p11_mult_21_n742) );
  XOR2_X2 p11_mult_21_U414 ( .A(reg2[10]), .B(p11_mult_21_n762), .Z(
        p11_mult_21_n725) );
  XOR2_X2 p11_mult_21_U413 ( .A(reg2[8]), .B(p11_mult_21_n760), .Z(
        p11_mult_21_n708) );
  XOR2_X2 p11_mult_21_U412 ( .A(reg2[6]), .B(p11_mult_21_n758), .Z(
        p11_mult_21_n691) );
  XOR2_X2 p11_mult_21_U411 ( .A(reg2[4]), .B(p11_mult_21_n771), .Z(
        p11_mult_21_n674) );
  INV_X1 p11_mult_21_U410 ( .A(reg2[0]), .ZN(p11_mult_21_n643) );
  INV_X1 p11_mult_21_U409 ( .A(p11_mult_21_n798), .ZN(p11_mult_21_n658) );
  HA_X1 p11_mult_21_U145 ( .A(p11_mult_21_n406), .B(p11_mult_21_n419), .CO(
        p11_mult_21_n315), .S(p11_mult_21_n316) );
  FA_X1 p11_mult_21_U144 ( .A(p11_mult_21_n418), .B(p11_mult_21_n393), .CI(
        p11_mult_21_n405), .CO(p11_mult_21_n313), .S(p11_mult_21_n314) );
  HA_X1 p11_mult_21_U143 ( .A(p11_mult_21_n321), .B(p11_mult_21_n392), .CO(
        p11_mult_21_n311), .S(p11_mult_21_n312) );
  FA_X1 p11_mult_21_U142 ( .A(p11_mult_21_n404), .B(p11_mult_21_n417), .CI(
        p11_mult_21_n312), .CO(p11_mult_21_n309), .S(p11_mult_21_n310) );
  FA_X1 p11_mult_21_U141 ( .A(p11_mult_21_n416), .B(p11_mult_21_n379), .CI(
        p11_mult_21_n403), .CO(p11_mult_21_n307), .S(p11_mult_21_n308) );
  FA_X1 p11_mult_21_U140 ( .A(p11_mult_21_n311), .B(p11_mult_21_n391), .CI(
        p11_mult_21_n308), .CO(p11_mult_21_n305), .S(p11_mult_21_n306) );
  HA_X1 p11_mult_21_U139 ( .A(p11_mult_21_n320), .B(p11_mult_21_n378), .CO(
        p11_mult_21_n303), .S(p11_mult_21_n304) );
  FA_X1 p11_mult_21_U138 ( .A(p11_mult_21_n390), .B(p11_mult_21_n415), .CI(
        p11_mult_21_n402), .CO(p11_mult_21_n301), .S(p11_mult_21_n302) );
  FA_X1 p11_mult_21_U137 ( .A(p11_mult_21_n307), .B(p11_mult_21_n304), .CI(
        p11_mult_21_n302), .CO(p11_mult_21_n299), .S(p11_mult_21_n300) );
  FA_X1 p11_mult_21_U136 ( .A(p11_mult_21_n389), .B(p11_mult_21_n365), .CI(
        p11_mult_21_n414), .CO(p11_mult_21_n297), .S(p11_mult_21_n298) );
  FA_X1 p11_mult_21_U135 ( .A(p11_mult_21_n377), .B(p11_mult_21_n401), .CI(
        p11_mult_21_n303), .CO(p11_mult_21_n295), .S(p11_mult_21_n296) );
  FA_X1 p11_mult_21_U134 ( .A(p11_mult_21_n298), .B(p11_mult_21_n301), .CI(
        p11_mult_21_n296), .CO(p11_mult_21_n293), .S(p11_mult_21_n294) );
  HA_X1 p11_mult_21_U133 ( .A(p11_mult_21_n319), .B(p11_mult_21_n364), .CO(
        p11_mult_21_n291), .S(p11_mult_21_n292) );
  FA_X1 p11_mult_21_U132 ( .A(p11_mult_21_n376), .B(p11_mult_21_n388), .CI(
        p11_mult_21_n400), .CO(p11_mult_21_n289), .S(p11_mult_21_n290) );
  FA_X1 p11_mult_21_U131 ( .A(p11_mult_21_n292), .B(p11_mult_21_n413), .CI(
        p11_mult_21_n297), .CO(p11_mult_21_n287), .S(p11_mult_21_n288) );
  FA_X1 p11_mult_21_U130 ( .A(p11_mult_21_n290), .B(p11_mult_21_n295), .CI(
        p11_mult_21_n288), .CO(p11_mult_21_n285), .S(p11_mult_21_n286) );
  FA_X1 p11_mult_21_U129 ( .A(p11_mult_21_n375), .B(p11_mult_21_n351), .CI(
        p11_mult_21_n412), .CO(p11_mult_21_n283), .S(p11_mult_21_n284) );
  FA_X1 p11_mult_21_U128 ( .A(p11_mult_21_n363), .B(p11_mult_21_n399), .CI(
        p11_mult_21_n387), .CO(p11_mult_21_n281), .S(p11_mult_21_n282) );
  FA_X1 p11_mult_21_U127 ( .A(p11_mult_21_n289), .B(p11_mult_21_n291), .CI(
        p11_mult_21_n284), .CO(p11_mult_21_n279), .S(p11_mult_21_n280) );
  FA_X1 p11_mult_21_U126 ( .A(p11_mult_21_n287), .B(p11_mult_21_n282), .CI(
        p11_mult_21_n280), .CO(p11_mult_21_n277), .S(p11_mult_21_n278) );
  HA_X1 p11_mult_21_U125 ( .A(p11_mult_21_n318), .B(p11_mult_21_n350), .CO(
        p11_mult_21_n275), .S(p11_mult_21_n276) );
  FA_X1 p11_mult_21_U124 ( .A(p11_mult_21_n362), .B(p11_mult_21_n386), .CI(
        p11_mult_21_n411), .CO(p11_mult_21_n273), .S(p11_mult_21_n274) );
  FA_X1 p11_mult_21_U123 ( .A(p11_mult_21_n374), .B(p11_mult_21_n398), .CI(
        p11_mult_21_n276), .CO(p11_mult_21_n271), .S(p11_mult_21_n272) );
  FA_X1 p11_mult_21_U122 ( .A(p11_mult_21_n281), .B(p11_mult_21_n283), .CI(
        p11_mult_21_n274), .CO(p11_mult_21_n269), .S(p11_mult_21_n270) );
  FA_X1 p11_mult_21_U121 ( .A(p11_mult_21_n279), .B(p11_mult_21_n272), .CI(
        p11_mult_21_n270), .CO(p11_mult_21_n267), .S(p11_mult_21_n268) );
  FA_X1 p11_mult_21_U120 ( .A(p11_mult_21_n361), .B(p11_mult_21_n337), .CI(
        p11_mult_21_n410), .CO(p11_mult_21_n265), .S(p11_mult_21_n266) );
  FA_X1 p11_mult_21_U109 ( .A(p11_mult_21_n349), .B(p11_mult_21_n397), .CI(
        p11_mult_21_n373), .CO(p11_mult_21_n263), .S(p11_mult_21_n264) );
  FA_X1 p11_mult_21_U108 ( .A(p11_mult_21_n275), .B(p11_mult_21_n385), .CI(
        p11_mult_21_n273), .CO(p11_mult_21_n261), .S(p11_mult_21_n262) );
  FA_X1 p11_mult_21_U107 ( .A(p11_mult_21_n264), .B(p11_mult_21_n266), .CI(
        p11_mult_21_n271), .CO(p11_mult_21_n259), .S(p11_mult_21_n260) );
  FA_X1 p11_mult_21_U106 ( .A(p11_mult_21_n262), .B(p11_mult_21_n269), .CI(
        p11_mult_21_n260), .CO(p11_mult_21_n257), .S(p11_mult_21_n258) );
  HA_X1 p11_mult_21_U105 ( .A(p11_mult_21_n317), .B(p11_mult_21_n336), .CO(
        p11_mult_21_n255), .S(p11_mult_21_n256) );
  FA_X1 p11_mult_21_U104 ( .A(p11_mult_21_n409), .B(p11_mult_21_n372), .CI(
        p11_mult_21_n396), .CO(p11_mult_21_n253), .S(p11_mult_21_n254) );
  FA_X1 p11_mult_21_U103 ( .A(p11_mult_21_n348), .B(p11_mult_21_n384), .CI(
        p11_mult_21_n360), .CO(p11_mult_21_n251), .S(p11_mult_21_n252) );
  FA_X1 p11_mult_21_U102 ( .A(p11_mult_21_n265), .B(p11_mult_21_n256), .CI(
        p11_mult_21_n263), .CO(p11_mult_21_n249), .S(p11_mult_21_n250) );
  FA_X1 p11_mult_21_U101 ( .A(p11_mult_21_n254), .B(p11_mult_21_n252), .CI(
        p11_mult_21_n261), .CO(p11_mult_21_n247), .S(p11_mult_21_n248) );
  FA_X1 p11_mult_21_U100 ( .A(p11_mult_21_n259), .B(p11_mult_21_n250), .CI(
        p11_mult_21_n248), .CO(p11_mult_21_n245), .S(p11_mult_21_n246) );
  FA_X1 p11_mult_21_U97 ( .A(p11_mult_21_n395), .B(p11_mult_21_n359), .CI(
        p11_mult_21_n408), .CO(p11_mult_21_n241), .S(p11_mult_21_n242) );
  FA_X1 p11_mult_21_U96 ( .A(p11_mult_21_n335), .B(p11_mult_21_n371), .CI(
        p11_mult_21_n255), .CO(p11_mult_21_n239), .S(p11_mult_21_n240) );
  FA_X1 p11_mult_21_U95 ( .A(p11_mult_21_n253), .B(p11_mult_21_n244), .CI(
        p11_mult_21_n251), .CO(p11_mult_21_n237), .S(p11_mult_21_n238) );
  FA_X1 p11_mult_21_U94 ( .A(p11_mult_21_n240), .B(p11_mult_21_n242), .CI(
        p11_mult_21_n249), .CO(p11_mult_21_n235), .S(p11_mult_21_n236) );
  FA_X1 p11_mult_21_U93 ( .A(p11_mult_21_n247), .B(p11_mult_21_n238), .CI(
        p11_mult_21_n236), .CO(p11_mult_21_n233), .S(p11_mult_21_n234) );
  FA_X1 p11_mult_21_U91 ( .A(p11_mult_21_n382), .B(p11_mult_21_n346), .CI(
        p11_mult_21_n232), .CO(p11_mult_21_n229), .S(p11_mult_21_n230) );
  FA_X1 p11_mult_21_U90 ( .A(p11_mult_21_n334), .B(p11_mult_21_n370), .CI(
        p11_mult_21_n358), .CO(p11_mult_21_n227), .S(p11_mult_21_n228) );
  FA_X1 p11_mult_21_U89 ( .A(p11_mult_21_n241), .B(p11_mult_21_n243), .CI(
        p11_mult_21_n239), .CO(p11_mult_21_n225), .S(p11_mult_21_n226) );
  FA_X1 p11_mult_21_U88 ( .A(p11_mult_21_n230), .B(p11_mult_21_n228), .CI(
        p11_mult_21_n237), .CO(p11_mult_21_n223), .S(p11_mult_21_n224) );
  FA_X1 p11_mult_21_U87 ( .A(p11_mult_21_n235), .B(p11_mult_21_n226), .CI(
        p11_mult_21_n224), .CO(p11_mult_21_n221), .S(p11_mult_21_n222) );
  FA_X1 p11_mult_21_U86 ( .A(p11_mult_21_n231), .B(p11_mult_21_n333), .CI(
        p11_mult_21_n394), .CO(p11_mult_21_n219), .S(p11_mult_21_n220) );
  FA_X1 p11_mult_21_U85 ( .A(p11_mult_21_n345), .B(p11_mult_21_n381), .CI(
        p11_mult_21_n357), .CO(p11_mult_21_n217), .S(p11_mult_21_n218) );
  FA_X1 p11_mult_21_U84 ( .A(p11_mult_21_n229), .B(p11_mult_21_n369), .CI(
        p11_mult_21_n227), .CO(p11_mult_21_n215), .S(p11_mult_21_n216) );
  FA_X1 p11_mult_21_U83 ( .A(p11_mult_21_n220), .B(p11_mult_21_n218), .CI(
        p11_mult_21_n225), .CO(p11_mult_21_n213), .S(p11_mult_21_n214) );
  FA_X1 p11_mult_21_U82 ( .A(p11_mult_21_n223), .B(p11_mult_21_n216), .CI(
        p11_mult_21_n214), .CO(p11_mult_21_n211), .S(p11_mult_21_n212) );
  FA_X1 p11_mult_21_U80 ( .A(p11_mult_21_n368), .B(p11_mult_21_n344), .CI(
        p11_mult_21_n210), .CO(p11_mult_21_n207), .S(p11_mult_21_n208) );
  FA_X1 p11_mult_21_U79 ( .A(p11_mult_21_n332), .B(p11_mult_21_n356), .CI(
        p11_mult_21_n219), .CO(p11_mult_21_n205), .S(p11_mult_21_n206) );
  FA_X1 p11_mult_21_U78 ( .A(p11_mult_21_n208), .B(p11_mult_21_n217), .CI(
        p11_mult_21_n215), .CO(p11_mult_21_n203), .S(p11_mult_21_n204) );
  FA_X1 p11_mult_21_U77 ( .A(p11_mult_21_n213), .B(p11_mult_21_n206), .CI(
        p11_mult_21_n204), .CO(p11_mult_21_n201), .S(p11_mult_21_n202) );
  FA_X1 p11_mult_21_U76 ( .A(p11_mult_21_n209), .B(p11_mult_21_n331), .CI(
        p11_mult_21_n380), .CO(p11_mult_21_n199), .S(p11_mult_21_n200) );
  FA_X1 p11_mult_21_U75 ( .A(p11_mult_21_n355), .B(p11_mult_21_n343), .CI(
        p11_mult_21_n367), .CO(p11_mult_21_n197), .S(p11_mult_21_n198) );
  FA_X1 p11_mult_21_U74 ( .A(p11_mult_21_n198), .B(p11_mult_21_n207), .CI(
        p11_mult_21_n200), .CO(p11_mult_21_n195), .S(p11_mult_21_n196) );
  FA_X1 p11_mult_21_U73 ( .A(p11_mult_21_n203), .B(p11_mult_21_n205), .CI(
        p11_mult_21_n196), .CO(p11_mult_21_n193), .S(p11_mult_21_n194) );
  FA_X1 p11_mult_21_U71 ( .A(p11_mult_21_n330), .B(p11_mult_21_n342), .CI(
        p11_mult_21_n192), .CO(p11_mult_21_n189), .S(p11_mult_21_n190) );
  FA_X1 p11_mult_21_U70 ( .A(p11_mult_21_n199), .B(p11_mult_21_n354), .CI(
        p11_mult_21_n197), .CO(p11_mult_21_n187), .S(p11_mult_21_n188) );
  FA_X1 p11_mult_21_U69 ( .A(p11_mult_21_n188), .B(p11_mult_21_n190), .CI(
        p11_mult_21_n195), .CO(p11_mult_21_n185), .S(p11_mult_21_n186) );
  FA_X1 p11_mult_21_U68 ( .A(p11_mult_21_n191), .B(p11_mult_21_n329), .CI(
        p11_mult_21_n366), .CO(p11_mult_21_n183), .S(p11_mult_21_n184) );
  FA_X1 p11_mult_21_U67 ( .A(p11_mult_21_n341), .B(p11_mult_21_n353), .CI(
        p11_mult_21_n189), .CO(p11_mult_21_n181), .S(p11_mult_21_n182) );
  FA_X1 p11_mult_21_U66 ( .A(p11_mult_21_n187), .B(p11_mult_21_n184), .CI(
        p11_mult_21_n182), .CO(p11_mult_21_n179), .S(p11_mult_21_n180) );
  FA_X1 p11_mult_21_U64 ( .A(p11_mult_21_n328), .B(p11_mult_21_n340), .CI(
        p11_mult_21_n178), .CO(p11_mult_21_n175), .S(p11_mult_21_n176) );
  FA_X1 p11_mult_21_U63 ( .A(p11_mult_21_n176), .B(p11_mult_21_n183), .CI(
        p11_mult_21_n181), .CO(p11_mult_21_n173), .S(p11_mult_21_n174) );
  FA_X1 p11_mult_21_U62 ( .A(p11_mult_21_n327), .B(p11_mult_21_n177), .CI(
        p11_mult_21_n352), .CO(p11_mult_21_n171), .S(p11_mult_21_n172) );
  FA_X1 p11_mult_21_U61 ( .A(p11_mult_21_n175), .B(p11_mult_21_n339), .CI(
        p11_mult_21_n172), .CO(p11_mult_21_n169), .S(p11_mult_21_n170) );
  FA_X1 p11_mult_21_U59 ( .A(p11_mult_21_n168), .B(p11_mult_21_n326), .CI(
        p11_mult_21_n171), .CO(p11_mult_21_n165), .S(p11_mult_21_n166) );
  FA_X1 p11_mult_21_U58 ( .A(p11_mult_21_n325), .B(p11_mult_21_n167), .CI(
        p11_mult_21_n338), .CO(p11_mult_21_n163), .S(p11_mult_21_n164) );
  FA_X1 p11_mult_21_U44 ( .A(p11_mult_21_n246), .B(p11_mult_21_n257), .CI(
        p11_mult_21_n149), .CO(p11_mult_21_n148), .S(temp6[0]) );
  FA_X1 p11_mult_21_U43 ( .A(p11_mult_21_n234), .B(p11_mult_21_n245), .CI(
        p11_mult_21_n148), .CO(p11_mult_21_n147), .S(temp6[1]) );
  FA_X1 p11_mult_21_U42 ( .A(p11_mult_21_n222), .B(p11_mult_21_n233), .CI(
        p11_mult_21_n147), .CO(p11_mult_21_n146), .S(temp6[2]) );
  FA_X1 p11_mult_21_U41 ( .A(p11_mult_21_n212), .B(p11_mult_21_n221), .CI(
        p11_mult_21_n146), .CO(p11_mult_21_n145), .S(temp6[3]) );
  FA_X1 p11_mult_21_U40 ( .A(p11_mult_21_n202), .B(p11_mult_21_n211), .CI(
        p11_mult_21_n145), .CO(p11_mult_21_n144), .S(temp6[4]) );
  FA_X1 p11_mult_21_U39 ( .A(p11_mult_21_n194), .B(p11_mult_21_n201), .CI(
        p11_mult_21_n144), .CO(p11_mult_21_n143), .S(temp6[5]) );
  FA_X1 p11_mult_21_U38 ( .A(p11_mult_21_n186), .B(p11_mult_21_n193), .CI(
        p11_mult_21_n143), .CO(p11_mult_21_n142), .S(temp6[6]) );
  FA_X1 p11_mult_21_U37 ( .A(p11_mult_21_n180), .B(p11_mult_21_n185), .CI(
        p11_mult_21_n142), .CO(p11_mult_21_n141), .S(temp6[7]) );
  FA_X1 p11_mult_21_U30 ( .A(p11_mult_21_n174), .B(p11_mult_21_n179), .CI(
        p11_mult_21_n141), .CO(p11_mult_21_n140), .S(temp6[8]) );
  FA_X1 p11_mult_21_U20 ( .A(p11_mult_21_n170), .B(p11_mult_21_n173), .CI(
        p11_mult_21_n140), .CO(p11_mult_21_n139), .S(temp6[9]) );
  FA_X1 p11_mult_21_U10 ( .A(p11_mult_21_n166), .B(p11_mult_21_n169), .CI(
        p11_mult_21_n139), .CO(p11_mult_21_n138), .S(temp6[10]) );
  FA_X1 p11_mult_21_U9 ( .A(p11_mult_21_n165), .B(p11_mult_21_n164), .CI(
        p11_mult_21_n138), .CO(p11_mult_21_n137), .S(temp6[11]) );
  FA_X1 p11_mult_21_U8 ( .A(p11_mult_21_n163), .B(p11_mult_21_n162), .CI(
        p11_mult_21_n137), .CO(p11_mult_21_n136), .S(temp6[12]) );
  XOR2_X1 p10_mult_21_U691 ( .A(reg4[2]), .B(reg4[1]), .Z(p10_mult_21_n798) );
  INV_X1 p10_mult_21_U690 ( .A(reg4[1]), .ZN(p10_mult_21_n655) );
  NOR2_X1 p10_mult_21_U689 ( .A1(p10_mult_21_n655), .A2(A2[1]), .ZN(
        p10_mult_21_n803) );
  INV_X1 p10_mult_21_U688 ( .A(p10_mult_21_n803), .ZN(p10_mult_21_n805) );
  NAND2_X1 p10_mult_21_U687 ( .A1(reg4[1]), .A2(p10_mult_21_n643), .ZN(
        p10_mult_21_n641) );
  XNOR2_X1 p10_mult_21_U686 ( .A(A2[2]), .B(reg4[1]), .ZN(p10_mult_21_n640) );
  OAI22_X1 p10_mult_21_U685 ( .A1(p10_mult_21_n805), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n640), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n804) );
  NAND2_X1 p10_mult_21_U684 ( .A1(p10_mult_21_n798), .A2(p10_mult_21_n804), 
        .ZN(p10_mult_21_n801) );
  NAND2_X1 p10_mult_21_U683 ( .A1(p10_mult_21_n803), .A2(p10_mult_21_n804), 
        .ZN(p10_mult_21_n802) );
  INV_X1 p10_mult_21_U682 ( .A(A2[0]), .ZN(p10_mult_21_n673) );
  MUX2_X1 p10_mult_21_U681 ( .A(p10_mult_21_n801), .B(p10_mult_21_n802), .S(
        p10_mult_21_n673), .Z(p10_mult_21_n800) );
  INV_X1 p10_mult_21_U680 ( .A(p10_mult_21_n800), .ZN(p10_mult_21_n795) );
  INV_X1 p10_mult_21_U679 ( .A(reg4[3]), .ZN(p10_mult_21_n771) );
  XNOR2_X1 p10_mult_21_U678 ( .A(p10_mult_21_n771), .B(reg4[2]), .ZN(
        p10_mult_21_n799) );
  NAND2_X1 p10_mult_21_U677 ( .A1(p10_mult_21_n658), .A2(p10_mult_21_n799), 
        .ZN(p10_mult_21_n657) );
  NAND3_X1 p10_mult_21_U676 ( .A1(p10_mult_21_n798), .A2(p10_mult_21_n673), 
        .A3(reg4[3]), .ZN(p10_mult_21_n797) );
  OAI21_X1 p10_mult_21_U675 ( .B1(p10_mult_21_n771), .B2(p10_mult_21_n657), 
        .A(p10_mult_21_n797), .ZN(p10_mult_21_n796) );
  AOI222_X1 p10_mult_21_U674 ( .A1(p10_mult_21_n795), .A2(p10_mult_21_n316), 
        .B1(p10_mult_21_n796), .B2(p10_mult_21_n795), .C1(p10_mult_21_n796), 
        .C2(p10_mult_21_n316), .ZN(p10_mult_21_n794) );
  INV_X1 p10_mult_21_U673 ( .A(p10_mult_21_n794), .ZN(p10_mult_21_n793) );
  AOI222_X1 p10_mult_21_U672 ( .A1(p10_mult_21_n793), .A2(p10_mult_21_n314), 
        .B1(p10_mult_21_n793), .B2(p10_mult_21_n315), .C1(p10_mult_21_n315), 
        .C2(p10_mult_21_n314), .ZN(p10_mult_21_n792) );
  INV_X1 p10_mult_21_U671 ( .A(p10_mult_21_n792), .ZN(p10_mult_21_n791) );
  AOI222_X1 p10_mult_21_U670 ( .A1(p10_mult_21_n791), .A2(p10_mult_21_n310), 
        .B1(p10_mult_21_n791), .B2(p10_mult_21_n313), .C1(p10_mult_21_n313), 
        .C2(p10_mult_21_n310), .ZN(p10_mult_21_n790) );
  INV_X1 p10_mult_21_U669 ( .A(p10_mult_21_n790), .ZN(p10_mult_21_n789) );
  AOI222_X1 p10_mult_21_U668 ( .A1(p10_mult_21_n789), .A2(p10_mult_21_n306), 
        .B1(p10_mult_21_n789), .B2(p10_mult_21_n309), .C1(p10_mult_21_n309), 
        .C2(p10_mult_21_n306), .ZN(p10_mult_21_n788) );
  INV_X1 p10_mult_21_U667 ( .A(p10_mult_21_n788), .ZN(p10_mult_21_n787) );
  AOI222_X1 p10_mult_21_U666 ( .A1(p10_mult_21_n787), .A2(p10_mult_21_n300), 
        .B1(p10_mult_21_n787), .B2(p10_mult_21_n305), .C1(p10_mult_21_n305), 
        .C2(p10_mult_21_n300), .ZN(p10_mult_21_n786) );
  INV_X1 p10_mult_21_U665 ( .A(p10_mult_21_n786), .ZN(p10_mult_21_n785) );
  AOI222_X1 p10_mult_21_U664 ( .A1(p10_mult_21_n785), .A2(p10_mult_21_n294), 
        .B1(p10_mult_21_n785), .B2(p10_mult_21_n299), .C1(p10_mult_21_n299), 
        .C2(p10_mult_21_n294), .ZN(p10_mult_21_n784) );
  INV_X1 p10_mult_21_U663 ( .A(p10_mult_21_n784), .ZN(p10_mult_21_n783) );
  AOI222_X1 p10_mult_21_U662 ( .A1(p10_mult_21_n783), .A2(p10_mult_21_n286), 
        .B1(p10_mult_21_n783), .B2(p10_mult_21_n293), .C1(p10_mult_21_n293), 
        .C2(p10_mult_21_n286), .ZN(p10_mult_21_n780) );
  INV_X1 p10_mult_21_U661 ( .A(p10_mult_21_n278), .ZN(p10_mult_21_n781) );
  INV_X1 p10_mult_21_U660 ( .A(p10_mult_21_n285), .ZN(p10_mult_21_n782) );
  OAI222_X1 p10_mult_21_U659 ( .A1(p10_mult_21_n780), .A2(p10_mult_21_n781), 
        .B1(p10_mult_21_n780), .B2(p10_mult_21_n782), .C1(p10_mult_21_n782), 
        .C2(p10_mult_21_n781), .ZN(p10_mult_21_n779) );
  AOI222_X1 p10_mult_21_U658 ( .A1(p10_mult_21_n779), .A2(p10_mult_21_n268), 
        .B1(p10_mult_21_n779), .B2(p10_mult_21_n277), .C1(p10_mult_21_n277), 
        .C2(p10_mult_21_n268), .ZN(p10_mult_21_n776) );
  INV_X1 p10_mult_21_U657 ( .A(p10_mult_21_n258), .ZN(p10_mult_21_n777) );
  INV_X1 p10_mult_21_U656 ( .A(p10_mult_21_n267), .ZN(p10_mult_21_n778) );
  OAI222_X1 p10_mult_21_U655 ( .A1(p10_mult_21_n776), .A2(p10_mult_21_n777), 
        .B1(p10_mult_21_n776), .B2(p10_mult_21_n778), .C1(p10_mult_21_n778), 
        .C2(p10_mult_21_n777), .ZN(p10_mult_21_n149) );
  XOR2_X1 p10_mult_21_U654 ( .A(A2[12]), .B(reg4[13]), .Z(p10_mult_21_n757) );
  INV_X1 p10_mult_21_U653 ( .A(reg4[11]), .ZN(p10_mult_21_n764) );
  INV_X1 p10_mult_21_U652 ( .A(reg4[13]), .ZN(p10_mult_21_n766) );
  XNOR2_X1 p10_mult_21_U651 ( .A(p10_mult_21_n766), .B(reg4[12]), .ZN(
        p10_mult_21_n775) );
  NAND2_X1 p10_mult_21_U650 ( .A1(p10_mult_21_n742), .A2(p10_mult_21_n775), 
        .ZN(p10_mult_21_n744) );
  INV_X1 p10_mult_21_U649 ( .A(p10_mult_21_n744), .ZN(p10_mult_21_n637) );
  INV_X1 p10_mult_21_U648 ( .A(p10_mult_21_n742), .ZN(p10_mult_21_n638) );
  XNOR2_X1 p10_mult_21_U647 ( .A(A2[13]), .B(p10_mult_21_n766), .ZN(
        p10_mult_21_n639) );
  AOI22_X1 p10_mult_21_U646 ( .A1(p10_mult_21_n757), .A2(p10_mult_21_n637), 
        .B1(p10_mult_21_n638), .B2(p10_mult_21_n639), .ZN(p10_mult_21_n162) );
  XNOR2_X1 p10_mult_21_U645 ( .A(A2[12]), .B(reg4[11]), .ZN(p10_mult_21_n739)
         );
  INV_X1 p10_mult_21_U644 ( .A(reg4[9]), .ZN(p10_mult_21_n762) );
  XNOR2_X1 p10_mult_21_U643 ( .A(p10_mult_21_n764), .B(reg4[10]), .ZN(
        p10_mult_21_n774) );
  NAND2_X1 p10_mult_21_U642 ( .A1(p10_mult_21_n725), .A2(p10_mult_21_n774), 
        .ZN(p10_mult_21_n727) );
  XNOR2_X1 p10_mult_21_U641 ( .A(A2[13]), .B(reg4[11]), .ZN(p10_mult_21_n741)
         );
  OAI22_X1 p10_mult_21_U640 ( .A1(p10_mult_21_n739), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n741), .ZN(p10_mult_21_n167) );
  INV_X1 p10_mult_21_U639 ( .A(p10_mult_21_n167), .ZN(p10_mult_21_n168) );
  XNOR2_X1 p10_mult_21_U638 ( .A(A2[12]), .B(reg4[9]), .ZN(p10_mult_21_n722)
         );
  INV_X1 p10_mult_21_U637 ( .A(reg4[7]), .ZN(p10_mult_21_n760) );
  XNOR2_X1 p10_mult_21_U636 ( .A(p10_mult_21_n762), .B(reg4[8]), .ZN(
        p10_mult_21_n773) );
  NAND2_X1 p10_mult_21_U635 ( .A1(p10_mult_21_n708), .A2(p10_mult_21_n773), 
        .ZN(p10_mult_21_n710) );
  XNOR2_X1 p10_mult_21_U634 ( .A(A2[13]), .B(reg4[9]), .ZN(p10_mult_21_n724)
         );
  OAI22_X1 p10_mult_21_U633 ( .A1(p10_mult_21_n722), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n724), .ZN(p10_mult_21_n177) );
  INV_X1 p10_mult_21_U632 ( .A(p10_mult_21_n177), .ZN(p10_mult_21_n178) );
  XNOR2_X1 p10_mult_21_U631 ( .A(A2[12]), .B(reg4[7]), .ZN(p10_mult_21_n705)
         );
  INV_X1 p10_mult_21_U630 ( .A(reg4[5]), .ZN(p10_mult_21_n758) );
  XNOR2_X1 p10_mult_21_U629 ( .A(p10_mult_21_n760), .B(reg4[6]), .ZN(
        p10_mult_21_n772) );
  NAND2_X1 p10_mult_21_U628 ( .A1(p10_mult_21_n691), .A2(p10_mult_21_n772), 
        .ZN(p10_mult_21_n693) );
  XNOR2_X1 p10_mult_21_U627 ( .A(A2[13]), .B(reg4[7]), .ZN(p10_mult_21_n707)
         );
  OAI22_X1 p10_mult_21_U626 ( .A1(p10_mult_21_n705), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n707), .ZN(p10_mult_21_n191) );
  INV_X1 p10_mult_21_U625 ( .A(p10_mult_21_n191), .ZN(p10_mult_21_n192) );
  XNOR2_X1 p10_mult_21_U624 ( .A(A2[12]), .B(reg4[5]), .ZN(p10_mult_21_n688)
         );
  XNOR2_X1 p10_mult_21_U623 ( .A(p10_mult_21_n758), .B(reg4[4]), .ZN(
        p10_mult_21_n770) );
  NAND2_X1 p10_mult_21_U622 ( .A1(p10_mult_21_n674), .A2(p10_mult_21_n770), 
        .ZN(p10_mult_21_n676) );
  XNOR2_X1 p10_mult_21_U621 ( .A(A2[13]), .B(reg4[5]), .ZN(p10_mult_21_n690)
         );
  OAI22_X1 p10_mult_21_U620 ( .A1(p10_mult_21_n688), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n690), .ZN(p10_mult_21_n209) );
  INV_X1 p10_mult_21_U619 ( .A(p10_mult_21_n209), .ZN(p10_mult_21_n210) );
  XNOR2_X1 p10_mult_21_U618 ( .A(A2[12]), .B(reg4[3]), .ZN(p10_mult_21_n670)
         );
  XNOR2_X1 p10_mult_21_U617 ( .A(A2[13]), .B(reg4[3]), .ZN(p10_mult_21_n672)
         );
  OAI22_X1 p10_mult_21_U616 ( .A1(p10_mult_21_n670), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n672), .ZN(p10_mult_21_n231) );
  INV_X1 p10_mult_21_U615 ( .A(p10_mult_21_n231), .ZN(p10_mult_21_n232) );
  XNOR2_X1 p10_mult_21_U614 ( .A(A2[3]), .B(reg4[11]), .ZN(p10_mult_21_n730)
         );
  XNOR2_X1 p10_mult_21_U613 ( .A(A2[4]), .B(reg4[11]), .ZN(p10_mult_21_n731)
         );
  OAI22_X1 p10_mult_21_U612 ( .A1(p10_mult_21_n730), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n731), .ZN(p10_mult_21_n768) );
  XNOR2_X1 p10_mult_21_U611 ( .A(A2[9]), .B(reg4[5]), .ZN(p10_mult_21_n685) );
  XNOR2_X1 p10_mult_21_U610 ( .A(A2[10]), .B(reg4[5]), .ZN(p10_mult_21_n686)
         );
  OAI22_X1 p10_mult_21_U609 ( .A1(p10_mult_21_n685), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n686), .ZN(p10_mult_21_n769) );
  OR2_X1 p10_mult_21_U608 ( .A1(p10_mult_21_n768), .A2(p10_mult_21_n769), .ZN(
        p10_mult_21_n243) );
  XNOR2_X1 p10_mult_21_U607 ( .A(p10_mult_21_n768), .B(p10_mult_21_n769), .ZN(
        p10_mult_21_n244) );
  NAND3_X1 p10_mult_21_U606 ( .A1(p10_mult_21_n638), .A2(p10_mult_21_n673), 
        .A3(reg4[13]), .ZN(p10_mult_21_n767) );
  OAI21_X1 p10_mult_21_U605 ( .B1(p10_mult_21_n766), .B2(p10_mult_21_n744), 
        .A(p10_mult_21_n767), .ZN(p10_mult_21_n317) );
  OR3_X1 p10_mult_21_U604 ( .A1(p10_mult_21_n725), .A2(A2[0]), .A3(
        p10_mult_21_n764), .ZN(p10_mult_21_n765) );
  OAI21_X1 p10_mult_21_U603 ( .B1(p10_mult_21_n764), .B2(p10_mult_21_n727), 
        .A(p10_mult_21_n765), .ZN(p10_mult_21_n318) );
  OR3_X1 p10_mult_21_U602 ( .A1(p10_mult_21_n708), .A2(A2[0]), .A3(
        p10_mult_21_n762), .ZN(p10_mult_21_n763) );
  OAI21_X1 p10_mult_21_U601 ( .B1(p10_mult_21_n762), .B2(p10_mult_21_n710), 
        .A(p10_mult_21_n763), .ZN(p10_mult_21_n319) );
  OR3_X1 p10_mult_21_U600 ( .A1(p10_mult_21_n691), .A2(A2[0]), .A3(
        p10_mult_21_n760), .ZN(p10_mult_21_n761) );
  OAI21_X1 p10_mult_21_U599 ( .B1(p10_mult_21_n760), .B2(p10_mult_21_n693), 
        .A(p10_mult_21_n761), .ZN(p10_mult_21_n320) );
  OR3_X1 p10_mult_21_U598 ( .A1(p10_mult_21_n674), .A2(A2[0]), .A3(
        p10_mult_21_n758), .ZN(p10_mult_21_n759) );
  OAI21_X1 p10_mult_21_U597 ( .B1(p10_mult_21_n758), .B2(p10_mult_21_n676), 
        .A(p10_mult_21_n759), .ZN(p10_mult_21_n321) );
  XNOR2_X1 p10_mult_21_U596 ( .A(A2[11]), .B(reg4[13]), .ZN(p10_mult_21_n755)
         );
  INV_X1 p10_mult_21_U595 ( .A(p10_mult_21_n757), .ZN(p10_mult_21_n756) );
  OAI22_X1 p10_mult_21_U594 ( .A1(p10_mult_21_n755), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n756), .ZN(p10_mult_21_n325) );
  XNOR2_X1 p10_mult_21_U593 ( .A(A2[10]), .B(reg4[13]), .ZN(p10_mult_21_n754)
         );
  OAI22_X1 p10_mult_21_U592 ( .A1(p10_mult_21_n754), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n755), .ZN(p10_mult_21_n326) );
  XNOR2_X1 p10_mult_21_U591 ( .A(A2[9]), .B(reg4[13]), .ZN(p10_mult_21_n753)
         );
  OAI22_X1 p10_mult_21_U590 ( .A1(p10_mult_21_n753), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n754), .ZN(p10_mult_21_n327) );
  XNOR2_X1 p10_mult_21_U589 ( .A(A2[8]), .B(reg4[13]), .ZN(p10_mult_21_n752)
         );
  OAI22_X1 p10_mult_21_U588 ( .A1(p10_mult_21_n752), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n753), .ZN(p10_mult_21_n328) );
  XNOR2_X1 p10_mult_21_U587 ( .A(A2[7]), .B(reg4[13]), .ZN(p10_mult_21_n751)
         );
  OAI22_X1 p10_mult_21_U586 ( .A1(p10_mult_21_n751), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n752), .ZN(p10_mult_21_n329) );
  XNOR2_X1 p10_mult_21_U585 ( .A(A2[6]), .B(reg4[13]), .ZN(p10_mult_21_n750)
         );
  OAI22_X1 p10_mult_21_U584 ( .A1(p10_mult_21_n750), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n751), .ZN(p10_mult_21_n330) );
  XNOR2_X1 p10_mult_21_U583 ( .A(A2[5]), .B(reg4[13]), .ZN(p10_mult_21_n749)
         );
  OAI22_X1 p10_mult_21_U582 ( .A1(p10_mult_21_n749), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n750), .ZN(p10_mult_21_n331) );
  XNOR2_X1 p10_mult_21_U581 ( .A(A2[4]), .B(reg4[13]), .ZN(p10_mult_21_n748)
         );
  OAI22_X1 p10_mult_21_U580 ( .A1(p10_mult_21_n748), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n749), .ZN(p10_mult_21_n332) );
  XNOR2_X1 p10_mult_21_U579 ( .A(A2[3]), .B(reg4[13]), .ZN(p10_mult_21_n747)
         );
  OAI22_X1 p10_mult_21_U578 ( .A1(p10_mult_21_n747), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n748), .ZN(p10_mult_21_n333) );
  XNOR2_X1 p10_mult_21_U577 ( .A(A2[2]), .B(reg4[13]), .ZN(p10_mult_21_n746)
         );
  OAI22_X1 p10_mult_21_U576 ( .A1(p10_mult_21_n746), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n747), .ZN(p10_mult_21_n334) );
  XNOR2_X1 p10_mult_21_U575 ( .A(A2[1]), .B(reg4[13]), .ZN(p10_mult_21_n745)
         );
  OAI22_X1 p10_mult_21_U574 ( .A1(p10_mult_21_n745), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n746), .ZN(p10_mult_21_n335) );
  XNOR2_X1 p10_mult_21_U573 ( .A(reg4[13]), .B(A2[0]), .ZN(p10_mult_21_n743)
         );
  OAI22_X1 p10_mult_21_U572 ( .A1(p10_mult_21_n743), .A2(p10_mult_21_n744), 
        .B1(p10_mult_21_n742), .B2(p10_mult_21_n745), .ZN(p10_mult_21_n336) );
  NOR2_X1 p10_mult_21_U571 ( .A1(p10_mult_21_n673), .A2(p10_mult_21_n742), 
        .ZN(p10_mult_21_n337) );
  AOI21_X1 p10_mult_21_U570 ( .B1(p10_mult_21_n727), .B2(p10_mult_21_n725), 
        .A(p10_mult_21_n741), .ZN(p10_mult_21_n740) );
  INV_X1 p10_mult_21_U569 ( .A(p10_mult_21_n740), .ZN(p10_mult_21_n338) );
  XNOR2_X1 p10_mult_21_U568 ( .A(A2[11]), .B(reg4[11]), .ZN(p10_mult_21_n738)
         );
  OAI22_X1 p10_mult_21_U567 ( .A1(p10_mult_21_n738), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n739), .ZN(p10_mult_21_n339) );
  XNOR2_X1 p10_mult_21_U566 ( .A(A2[10]), .B(reg4[11]), .ZN(p10_mult_21_n737)
         );
  OAI22_X1 p10_mult_21_U565 ( .A1(p10_mult_21_n737), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n738), .ZN(p10_mult_21_n340) );
  XNOR2_X1 p10_mult_21_U564 ( .A(A2[9]), .B(reg4[11]), .ZN(p10_mult_21_n736)
         );
  OAI22_X1 p10_mult_21_U563 ( .A1(p10_mult_21_n736), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n737), .ZN(p10_mult_21_n341) );
  XNOR2_X1 p10_mult_21_U562 ( .A(A2[8]), .B(reg4[11]), .ZN(p10_mult_21_n735)
         );
  OAI22_X1 p10_mult_21_U561 ( .A1(p10_mult_21_n735), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n736), .ZN(p10_mult_21_n342) );
  XNOR2_X1 p10_mult_21_U560 ( .A(A2[7]), .B(reg4[11]), .ZN(p10_mult_21_n734)
         );
  OAI22_X1 p10_mult_21_U559 ( .A1(p10_mult_21_n734), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n735), .ZN(p10_mult_21_n343) );
  XNOR2_X1 p10_mult_21_U558 ( .A(A2[6]), .B(reg4[11]), .ZN(p10_mult_21_n733)
         );
  OAI22_X1 p10_mult_21_U557 ( .A1(p10_mult_21_n733), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n734), .ZN(p10_mult_21_n344) );
  XNOR2_X1 p10_mult_21_U556 ( .A(A2[5]), .B(reg4[11]), .ZN(p10_mult_21_n732)
         );
  OAI22_X1 p10_mult_21_U555 ( .A1(p10_mult_21_n732), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n733), .ZN(p10_mult_21_n345) );
  OAI22_X1 p10_mult_21_U554 ( .A1(p10_mult_21_n731), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n732), .ZN(p10_mult_21_n346) );
  XNOR2_X1 p10_mult_21_U553 ( .A(A2[2]), .B(reg4[11]), .ZN(p10_mult_21_n729)
         );
  OAI22_X1 p10_mult_21_U552 ( .A1(p10_mult_21_n729), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n730), .ZN(p10_mult_21_n348) );
  XNOR2_X1 p10_mult_21_U551 ( .A(A2[1]), .B(reg4[11]), .ZN(p10_mult_21_n728)
         );
  OAI22_X1 p10_mult_21_U550 ( .A1(p10_mult_21_n728), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n729), .ZN(p10_mult_21_n349) );
  XNOR2_X1 p10_mult_21_U549 ( .A(reg4[11]), .B(A2[0]), .ZN(p10_mult_21_n726)
         );
  OAI22_X1 p10_mult_21_U548 ( .A1(p10_mult_21_n726), .A2(p10_mult_21_n727), 
        .B1(p10_mult_21_n725), .B2(p10_mult_21_n728), .ZN(p10_mult_21_n350) );
  NOR2_X1 p10_mult_21_U547 ( .A1(p10_mult_21_n673), .A2(p10_mult_21_n725), 
        .ZN(p10_mult_21_n351) );
  AOI21_X1 p10_mult_21_U546 ( .B1(p10_mult_21_n710), .B2(p10_mult_21_n708), 
        .A(p10_mult_21_n724), .ZN(p10_mult_21_n723) );
  INV_X1 p10_mult_21_U545 ( .A(p10_mult_21_n723), .ZN(p10_mult_21_n352) );
  XNOR2_X1 p10_mult_21_U544 ( .A(A2[11]), .B(reg4[9]), .ZN(p10_mult_21_n721)
         );
  OAI22_X1 p10_mult_21_U543 ( .A1(p10_mult_21_n721), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n722), .ZN(p10_mult_21_n353) );
  XNOR2_X1 p10_mult_21_U542 ( .A(A2[10]), .B(reg4[9]), .ZN(p10_mult_21_n720)
         );
  OAI22_X1 p10_mult_21_U541 ( .A1(p10_mult_21_n720), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n721), .ZN(p10_mult_21_n354) );
  XNOR2_X1 p10_mult_21_U540 ( .A(A2[9]), .B(reg4[9]), .ZN(p10_mult_21_n719) );
  OAI22_X1 p10_mult_21_U539 ( .A1(p10_mult_21_n719), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n720), .ZN(p10_mult_21_n355) );
  XNOR2_X1 p10_mult_21_U538 ( .A(A2[8]), .B(reg4[9]), .ZN(p10_mult_21_n718) );
  OAI22_X1 p10_mult_21_U537 ( .A1(p10_mult_21_n718), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n719), .ZN(p10_mult_21_n356) );
  XNOR2_X1 p10_mult_21_U536 ( .A(A2[7]), .B(reg4[9]), .ZN(p10_mult_21_n717) );
  OAI22_X1 p10_mult_21_U535 ( .A1(p10_mult_21_n717), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n718), .ZN(p10_mult_21_n357) );
  XNOR2_X1 p10_mult_21_U534 ( .A(A2[6]), .B(reg4[9]), .ZN(p10_mult_21_n716) );
  OAI22_X1 p10_mult_21_U533 ( .A1(p10_mult_21_n716), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n717), .ZN(p10_mult_21_n358) );
  XNOR2_X1 p10_mult_21_U532 ( .A(A2[5]), .B(reg4[9]), .ZN(p10_mult_21_n715) );
  OAI22_X1 p10_mult_21_U531 ( .A1(p10_mult_21_n715), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n716), .ZN(p10_mult_21_n359) );
  XNOR2_X1 p10_mult_21_U530 ( .A(A2[4]), .B(reg4[9]), .ZN(p10_mult_21_n714) );
  OAI22_X1 p10_mult_21_U529 ( .A1(p10_mult_21_n714), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n715), .ZN(p10_mult_21_n360) );
  XNOR2_X1 p10_mult_21_U528 ( .A(A2[3]), .B(reg4[9]), .ZN(p10_mult_21_n713) );
  OAI22_X1 p10_mult_21_U527 ( .A1(p10_mult_21_n713), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n714), .ZN(p10_mult_21_n361) );
  XNOR2_X1 p10_mult_21_U526 ( .A(A2[2]), .B(reg4[9]), .ZN(p10_mult_21_n712) );
  OAI22_X1 p10_mult_21_U525 ( .A1(p10_mult_21_n712), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n713), .ZN(p10_mult_21_n362) );
  XNOR2_X1 p10_mult_21_U524 ( .A(A2[1]), .B(reg4[9]), .ZN(p10_mult_21_n711) );
  OAI22_X1 p10_mult_21_U523 ( .A1(p10_mult_21_n711), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n712), .ZN(p10_mult_21_n363) );
  XNOR2_X1 p10_mult_21_U522 ( .A(reg4[9]), .B(A2[0]), .ZN(p10_mult_21_n709) );
  OAI22_X1 p10_mult_21_U521 ( .A1(p10_mult_21_n709), .A2(p10_mult_21_n710), 
        .B1(p10_mult_21_n708), .B2(p10_mult_21_n711), .ZN(p10_mult_21_n364) );
  NOR2_X1 p10_mult_21_U520 ( .A1(p10_mult_21_n673), .A2(p10_mult_21_n708), 
        .ZN(p10_mult_21_n365) );
  AOI21_X1 p10_mult_21_U519 ( .B1(p10_mult_21_n693), .B2(p10_mult_21_n691), 
        .A(p10_mult_21_n707), .ZN(p10_mult_21_n706) );
  INV_X1 p10_mult_21_U518 ( .A(p10_mult_21_n706), .ZN(p10_mult_21_n366) );
  XNOR2_X1 p10_mult_21_U517 ( .A(A2[11]), .B(reg4[7]), .ZN(p10_mult_21_n704)
         );
  OAI22_X1 p10_mult_21_U516 ( .A1(p10_mult_21_n704), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n705), .ZN(p10_mult_21_n367) );
  XNOR2_X1 p10_mult_21_U515 ( .A(A2[10]), .B(reg4[7]), .ZN(p10_mult_21_n703)
         );
  OAI22_X1 p10_mult_21_U514 ( .A1(p10_mult_21_n703), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n704), .ZN(p10_mult_21_n368) );
  XNOR2_X1 p10_mult_21_U513 ( .A(A2[9]), .B(reg4[7]), .ZN(p10_mult_21_n702) );
  OAI22_X1 p10_mult_21_U512 ( .A1(p10_mult_21_n702), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n703), .ZN(p10_mult_21_n369) );
  XNOR2_X1 p10_mult_21_U511 ( .A(A2[8]), .B(reg4[7]), .ZN(p10_mult_21_n701) );
  OAI22_X1 p10_mult_21_U510 ( .A1(p10_mult_21_n701), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n702), .ZN(p10_mult_21_n370) );
  XNOR2_X1 p10_mult_21_U509 ( .A(A2[7]), .B(reg4[7]), .ZN(p10_mult_21_n700) );
  OAI22_X1 p10_mult_21_U508 ( .A1(p10_mult_21_n700), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n701), .ZN(p10_mult_21_n371) );
  XNOR2_X1 p10_mult_21_U507 ( .A(A2[6]), .B(reg4[7]), .ZN(p10_mult_21_n699) );
  OAI22_X1 p10_mult_21_U506 ( .A1(p10_mult_21_n699), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n700), .ZN(p10_mult_21_n372) );
  XNOR2_X1 p10_mult_21_U505 ( .A(A2[5]), .B(reg4[7]), .ZN(p10_mult_21_n698) );
  OAI22_X1 p10_mult_21_U504 ( .A1(p10_mult_21_n698), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n699), .ZN(p10_mult_21_n373) );
  XNOR2_X1 p10_mult_21_U503 ( .A(A2[4]), .B(reg4[7]), .ZN(p10_mult_21_n697) );
  OAI22_X1 p10_mult_21_U502 ( .A1(p10_mult_21_n697), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n698), .ZN(p10_mult_21_n374) );
  XNOR2_X1 p10_mult_21_U501 ( .A(A2[3]), .B(reg4[7]), .ZN(p10_mult_21_n696) );
  OAI22_X1 p10_mult_21_U500 ( .A1(p10_mult_21_n696), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n697), .ZN(p10_mult_21_n375) );
  XNOR2_X1 p10_mult_21_U499 ( .A(A2[2]), .B(reg4[7]), .ZN(p10_mult_21_n695) );
  OAI22_X1 p10_mult_21_U498 ( .A1(p10_mult_21_n695), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n696), .ZN(p10_mult_21_n376) );
  XNOR2_X1 p10_mult_21_U497 ( .A(A2[1]), .B(reg4[7]), .ZN(p10_mult_21_n694) );
  OAI22_X1 p10_mult_21_U496 ( .A1(p10_mult_21_n694), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n695), .ZN(p10_mult_21_n377) );
  XNOR2_X1 p10_mult_21_U495 ( .A(reg4[7]), .B(A2[0]), .ZN(p10_mult_21_n692) );
  OAI22_X1 p10_mult_21_U494 ( .A1(p10_mult_21_n692), .A2(p10_mult_21_n693), 
        .B1(p10_mult_21_n691), .B2(p10_mult_21_n694), .ZN(p10_mult_21_n378) );
  NOR2_X1 p10_mult_21_U493 ( .A1(p10_mult_21_n673), .A2(p10_mult_21_n691), 
        .ZN(p10_mult_21_n379) );
  AOI21_X1 p10_mult_21_U492 ( .B1(p10_mult_21_n676), .B2(p10_mult_21_n674), 
        .A(p10_mult_21_n690), .ZN(p10_mult_21_n689) );
  INV_X1 p10_mult_21_U491 ( .A(p10_mult_21_n689), .ZN(p10_mult_21_n380) );
  XNOR2_X1 p10_mult_21_U490 ( .A(A2[11]), .B(reg4[5]), .ZN(p10_mult_21_n687)
         );
  OAI22_X1 p10_mult_21_U489 ( .A1(p10_mult_21_n687), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n688), .ZN(p10_mult_21_n381) );
  OAI22_X1 p10_mult_21_U488 ( .A1(p10_mult_21_n686), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n687), .ZN(p10_mult_21_n382) );
  XNOR2_X1 p10_mult_21_U487 ( .A(A2[8]), .B(reg4[5]), .ZN(p10_mult_21_n684) );
  OAI22_X1 p10_mult_21_U486 ( .A1(p10_mult_21_n684), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n685), .ZN(p10_mult_21_n384) );
  XNOR2_X1 p10_mult_21_U485 ( .A(A2[7]), .B(reg4[5]), .ZN(p10_mult_21_n683) );
  OAI22_X1 p10_mult_21_U484 ( .A1(p10_mult_21_n683), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n684), .ZN(p10_mult_21_n385) );
  XNOR2_X1 p10_mult_21_U483 ( .A(A2[6]), .B(reg4[5]), .ZN(p10_mult_21_n682) );
  OAI22_X1 p10_mult_21_U482 ( .A1(p10_mult_21_n682), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n683), .ZN(p10_mult_21_n386) );
  XNOR2_X1 p10_mult_21_U481 ( .A(A2[5]), .B(reg4[5]), .ZN(p10_mult_21_n681) );
  OAI22_X1 p10_mult_21_U480 ( .A1(p10_mult_21_n681), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n682), .ZN(p10_mult_21_n387) );
  XNOR2_X1 p10_mult_21_U479 ( .A(A2[4]), .B(reg4[5]), .ZN(p10_mult_21_n680) );
  OAI22_X1 p10_mult_21_U478 ( .A1(p10_mult_21_n680), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n681), .ZN(p10_mult_21_n388) );
  XNOR2_X1 p10_mult_21_U477 ( .A(A2[3]), .B(reg4[5]), .ZN(p10_mult_21_n679) );
  OAI22_X1 p10_mult_21_U476 ( .A1(p10_mult_21_n679), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n680), .ZN(p10_mult_21_n389) );
  XNOR2_X1 p10_mult_21_U475 ( .A(A2[2]), .B(reg4[5]), .ZN(p10_mult_21_n678) );
  OAI22_X1 p10_mult_21_U474 ( .A1(p10_mult_21_n678), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n679), .ZN(p10_mult_21_n390) );
  XNOR2_X1 p10_mult_21_U473 ( .A(A2[1]), .B(reg4[5]), .ZN(p10_mult_21_n677) );
  OAI22_X1 p10_mult_21_U472 ( .A1(p10_mult_21_n677), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n678), .ZN(p10_mult_21_n391) );
  XNOR2_X1 p10_mult_21_U471 ( .A(reg4[5]), .B(A2[0]), .ZN(p10_mult_21_n675) );
  OAI22_X1 p10_mult_21_U470 ( .A1(p10_mult_21_n675), .A2(p10_mult_21_n676), 
        .B1(p10_mult_21_n674), .B2(p10_mult_21_n677), .ZN(p10_mult_21_n392) );
  NOR2_X1 p10_mult_21_U469 ( .A1(p10_mult_21_n673), .A2(p10_mult_21_n674), 
        .ZN(p10_mult_21_n393) );
  AOI21_X1 p10_mult_21_U468 ( .B1(p10_mult_21_n657), .B2(p10_mult_21_n658), 
        .A(p10_mult_21_n672), .ZN(p10_mult_21_n671) );
  INV_X1 p10_mult_21_U467 ( .A(p10_mult_21_n671), .ZN(p10_mult_21_n394) );
  XNOR2_X1 p10_mult_21_U466 ( .A(A2[11]), .B(reg4[3]), .ZN(p10_mult_21_n669)
         );
  OAI22_X1 p10_mult_21_U465 ( .A1(p10_mult_21_n669), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n670), .ZN(p10_mult_21_n395) );
  XNOR2_X1 p10_mult_21_U464 ( .A(A2[10]), .B(reg4[3]), .ZN(p10_mult_21_n668)
         );
  OAI22_X1 p10_mult_21_U463 ( .A1(p10_mult_21_n668), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n669), .ZN(p10_mult_21_n396) );
  XNOR2_X1 p10_mult_21_U462 ( .A(A2[9]), .B(reg4[3]), .ZN(p10_mult_21_n667) );
  OAI22_X1 p10_mult_21_U461 ( .A1(p10_mult_21_n667), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n668), .ZN(p10_mult_21_n397) );
  XNOR2_X1 p10_mult_21_U460 ( .A(A2[8]), .B(reg4[3]), .ZN(p10_mult_21_n666) );
  OAI22_X1 p10_mult_21_U459 ( .A1(p10_mult_21_n666), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n667), .ZN(p10_mult_21_n398) );
  XNOR2_X1 p10_mult_21_U458 ( .A(A2[7]), .B(reg4[3]), .ZN(p10_mult_21_n665) );
  OAI22_X1 p10_mult_21_U457 ( .A1(p10_mult_21_n665), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n666), .ZN(p10_mult_21_n399) );
  XNOR2_X1 p10_mult_21_U456 ( .A(A2[6]), .B(reg4[3]), .ZN(p10_mult_21_n664) );
  OAI22_X1 p10_mult_21_U455 ( .A1(p10_mult_21_n664), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n665), .ZN(p10_mult_21_n400) );
  XNOR2_X1 p10_mult_21_U454 ( .A(A2[5]), .B(reg4[3]), .ZN(p10_mult_21_n663) );
  OAI22_X1 p10_mult_21_U453 ( .A1(p10_mult_21_n663), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n664), .ZN(p10_mult_21_n401) );
  XNOR2_X1 p10_mult_21_U452 ( .A(A2[4]), .B(reg4[3]), .ZN(p10_mult_21_n662) );
  OAI22_X1 p10_mult_21_U451 ( .A1(p10_mult_21_n662), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n663), .ZN(p10_mult_21_n402) );
  XNOR2_X1 p10_mult_21_U450 ( .A(A2[3]), .B(reg4[3]), .ZN(p10_mult_21_n661) );
  OAI22_X1 p10_mult_21_U449 ( .A1(p10_mult_21_n661), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n662), .ZN(p10_mult_21_n403) );
  XNOR2_X1 p10_mult_21_U448 ( .A(A2[2]), .B(reg4[3]), .ZN(p10_mult_21_n660) );
  OAI22_X1 p10_mult_21_U447 ( .A1(p10_mult_21_n660), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n661), .ZN(p10_mult_21_n404) );
  XNOR2_X1 p10_mult_21_U446 ( .A(A2[1]), .B(reg4[3]), .ZN(p10_mult_21_n659) );
  OAI22_X1 p10_mult_21_U445 ( .A1(p10_mult_21_n659), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n660), .ZN(p10_mult_21_n405) );
  XNOR2_X1 p10_mult_21_U444 ( .A(reg4[3]), .B(A2[0]), .ZN(p10_mult_21_n656) );
  OAI22_X1 p10_mult_21_U443 ( .A1(p10_mult_21_n656), .A2(p10_mult_21_n657), 
        .B1(p10_mult_21_n658), .B2(p10_mult_21_n659), .ZN(p10_mult_21_n406) );
  XOR2_X1 p10_mult_21_U442 ( .A(A2[13]), .B(p10_mult_21_n655), .Z(
        p10_mult_21_n653) );
  AOI21_X1 p10_mult_21_U441 ( .B1(p10_mult_21_n641), .B2(p10_mult_21_n643), 
        .A(p10_mult_21_n653), .ZN(p10_mult_21_n654) );
  INV_X1 p10_mult_21_U440 ( .A(p10_mult_21_n654), .ZN(p10_mult_21_n408) );
  XNOR2_X1 p10_mult_21_U439 ( .A(A2[12]), .B(reg4[1]), .ZN(p10_mult_21_n652)
         );
  OAI22_X1 p10_mult_21_U438 ( .A1(p10_mult_21_n652), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n653), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n409) );
  XNOR2_X1 p10_mult_21_U437 ( .A(A2[11]), .B(reg4[1]), .ZN(p10_mult_21_n651)
         );
  OAI22_X1 p10_mult_21_U436 ( .A1(p10_mult_21_n651), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n652), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n410) );
  XNOR2_X1 p10_mult_21_U435 ( .A(A2[10]), .B(reg4[1]), .ZN(p10_mult_21_n650)
         );
  OAI22_X1 p10_mult_21_U434 ( .A1(p10_mult_21_n650), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n651), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n411) );
  XNOR2_X1 p10_mult_21_U433 ( .A(A2[9]), .B(reg4[1]), .ZN(p10_mult_21_n649) );
  OAI22_X1 p10_mult_21_U432 ( .A1(p10_mult_21_n649), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n650), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n412) );
  XNOR2_X1 p10_mult_21_U431 ( .A(A2[8]), .B(reg4[1]), .ZN(p10_mult_21_n648) );
  OAI22_X1 p10_mult_21_U430 ( .A1(p10_mult_21_n648), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n649), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n413) );
  XNOR2_X1 p10_mult_21_U429 ( .A(A2[7]), .B(reg4[1]), .ZN(p10_mult_21_n647) );
  OAI22_X1 p10_mult_21_U428 ( .A1(p10_mult_21_n647), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n648), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n414) );
  XNOR2_X1 p10_mult_21_U427 ( .A(A2[6]), .B(reg4[1]), .ZN(p10_mult_21_n646) );
  OAI22_X1 p10_mult_21_U426 ( .A1(p10_mult_21_n646), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n647), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n415) );
  XNOR2_X1 p10_mult_21_U425 ( .A(A2[5]), .B(reg4[1]), .ZN(p10_mult_21_n645) );
  OAI22_X1 p10_mult_21_U424 ( .A1(p10_mult_21_n645), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n646), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n416) );
  XNOR2_X1 p10_mult_21_U423 ( .A(A2[4]), .B(reg4[1]), .ZN(p10_mult_21_n644) );
  OAI22_X1 p10_mult_21_U422 ( .A1(p10_mult_21_n644), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n645), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n417) );
  XNOR2_X1 p10_mult_21_U421 ( .A(A2[3]), .B(reg4[1]), .ZN(p10_mult_21_n642) );
  OAI22_X1 p10_mult_21_U420 ( .A1(p10_mult_21_n642), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n644), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n418) );
  OAI22_X1 p10_mult_21_U419 ( .A1(p10_mult_21_n640), .A2(p10_mult_21_n641), 
        .B1(p10_mult_21_n642), .B2(p10_mult_21_n643), .ZN(p10_mult_21_n419) );
  OAI21_X1 p10_mult_21_U418 ( .B1(p10_mult_21_n637), .B2(p10_mult_21_n638), 
        .A(p10_mult_21_n639), .ZN(p10_mult_21_n636) );
  XOR2_X1 p10_mult_21_U417 ( .A(p10_mult_21_n636), .B(p10_mult_21_n136), .Z(
        p10_mult_21_n635) );
  XNOR2_X1 p10_mult_21_U416 ( .A(p10_mult_21_n162), .B(p10_mult_21_n635), .ZN(
        temp5[13]) );
  XOR2_X2 p10_mult_21_U415 ( .A(reg4[12]), .B(p10_mult_21_n764), .Z(
        p10_mult_21_n742) );
  XOR2_X2 p10_mult_21_U414 ( .A(reg4[10]), .B(p10_mult_21_n762), .Z(
        p10_mult_21_n725) );
  XOR2_X2 p10_mult_21_U413 ( .A(reg4[8]), .B(p10_mult_21_n760), .Z(
        p10_mult_21_n708) );
  XOR2_X2 p10_mult_21_U412 ( .A(reg4[6]), .B(p10_mult_21_n758), .Z(
        p10_mult_21_n691) );
  XOR2_X2 p10_mult_21_U411 ( .A(reg4[4]), .B(p10_mult_21_n771), .Z(
        p10_mult_21_n674) );
  INV_X1 p10_mult_21_U410 ( .A(reg4[0]), .ZN(p10_mult_21_n643) );
  INV_X1 p10_mult_21_U409 ( .A(p10_mult_21_n798), .ZN(p10_mult_21_n658) );
  HA_X1 p10_mult_21_U145 ( .A(p10_mult_21_n406), .B(p10_mult_21_n419), .CO(
        p10_mult_21_n315), .S(p10_mult_21_n316) );
  FA_X1 p10_mult_21_U144 ( .A(p10_mult_21_n418), .B(p10_mult_21_n393), .CI(
        p10_mult_21_n405), .CO(p10_mult_21_n313), .S(p10_mult_21_n314) );
  HA_X1 p10_mult_21_U143 ( .A(p10_mult_21_n321), .B(p10_mult_21_n392), .CO(
        p10_mult_21_n311), .S(p10_mult_21_n312) );
  FA_X1 p10_mult_21_U142 ( .A(p10_mult_21_n404), .B(p10_mult_21_n417), .CI(
        p10_mult_21_n312), .CO(p10_mult_21_n309), .S(p10_mult_21_n310) );
  FA_X1 p10_mult_21_U141 ( .A(p10_mult_21_n416), .B(p10_mult_21_n379), .CI(
        p10_mult_21_n403), .CO(p10_mult_21_n307), .S(p10_mult_21_n308) );
  FA_X1 p10_mult_21_U140 ( .A(p10_mult_21_n311), .B(p10_mult_21_n391), .CI(
        p10_mult_21_n308), .CO(p10_mult_21_n305), .S(p10_mult_21_n306) );
  HA_X1 p10_mult_21_U139 ( .A(p10_mult_21_n320), .B(p10_mult_21_n378), .CO(
        p10_mult_21_n303), .S(p10_mult_21_n304) );
  FA_X1 p10_mult_21_U138 ( .A(p10_mult_21_n390), .B(p10_mult_21_n415), .CI(
        p10_mult_21_n402), .CO(p10_mult_21_n301), .S(p10_mult_21_n302) );
  FA_X1 p10_mult_21_U137 ( .A(p10_mult_21_n307), .B(p10_mult_21_n304), .CI(
        p10_mult_21_n302), .CO(p10_mult_21_n299), .S(p10_mult_21_n300) );
  FA_X1 p10_mult_21_U136 ( .A(p10_mult_21_n389), .B(p10_mult_21_n365), .CI(
        p10_mult_21_n414), .CO(p10_mult_21_n297), .S(p10_mult_21_n298) );
  FA_X1 p10_mult_21_U135 ( .A(p10_mult_21_n377), .B(p10_mult_21_n401), .CI(
        p10_mult_21_n303), .CO(p10_mult_21_n295), .S(p10_mult_21_n296) );
  FA_X1 p10_mult_21_U134 ( .A(p10_mult_21_n298), .B(p10_mult_21_n301), .CI(
        p10_mult_21_n296), .CO(p10_mult_21_n293), .S(p10_mult_21_n294) );
  HA_X1 p10_mult_21_U133 ( .A(p10_mult_21_n319), .B(p10_mult_21_n364), .CO(
        p10_mult_21_n291), .S(p10_mult_21_n292) );
  FA_X1 p10_mult_21_U132 ( .A(p10_mult_21_n376), .B(p10_mult_21_n388), .CI(
        p10_mult_21_n400), .CO(p10_mult_21_n289), .S(p10_mult_21_n290) );
  FA_X1 p10_mult_21_U131 ( .A(p10_mult_21_n292), .B(p10_mult_21_n413), .CI(
        p10_mult_21_n297), .CO(p10_mult_21_n287), .S(p10_mult_21_n288) );
  FA_X1 p10_mult_21_U130 ( .A(p10_mult_21_n290), .B(p10_mult_21_n295), .CI(
        p10_mult_21_n288), .CO(p10_mult_21_n285), .S(p10_mult_21_n286) );
  FA_X1 p10_mult_21_U129 ( .A(p10_mult_21_n375), .B(p10_mult_21_n351), .CI(
        p10_mult_21_n412), .CO(p10_mult_21_n283), .S(p10_mult_21_n284) );
  FA_X1 p10_mult_21_U128 ( .A(p10_mult_21_n363), .B(p10_mult_21_n399), .CI(
        p10_mult_21_n387), .CO(p10_mult_21_n281), .S(p10_mult_21_n282) );
  FA_X1 p10_mult_21_U127 ( .A(p10_mult_21_n289), .B(p10_mult_21_n291), .CI(
        p10_mult_21_n284), .CO(p10_mult_21_n279), .S(p10_mult_21_n280) );
  FA_X1 p10_mult_21_U126 ( .A(p10_mult_21_n287), .B(p10_mult_21_n282), .CI(
        p10_mult_21_n280), .CO(p10_mult_21_n277), .S(p10_mult_21_n278) );
  HA_X1 p10_mult_21_U125 ( .A(p10_mult_21_n318), .B(p10_mult_21_n350), .CO(
        p10_mult_21_n275), .S(p10_mult_21_n276) );
  FA_X1 p10_mult_21_U124 ( .A(p10_mult_21_n362), .B(p10_mult_21_n386), .CI(
        p10_mult_21_n411), .CO(p10_mult_21_n273), .S(p10_mult_21_n274) );
  FA_X1 p10_mult_21_U123 ( .A(p10_mult_21_n374), .B(p10_mult_21_n398), .CI(
        p10_mult_21_n276), .CO(p10_mult_21_n271), .S(p10_mult_21_n272) );
  FA_X1 p10_mult_21_U122 ( .A(p10_mult_21_n281), .B(p10_mult_21_n283), .CI(
        p10_mult_21_n274), .CO(p10_mult_21_n269), .S(p10_mult_21_n270) );
  FA_X1 p10_mult_21_U121 ( .A(p10_mult_21_n279), .B(p10_mult_21_n272), .CI(
        p10_mult_21_n270), .CO(p10_mult_21_n267), .S(p10_mult_21_n268) );
  FA_X1 p10_mult_21_U120 ( .A(p10_mult_21_n361), .B(p10_mult_21_n337), .CI(
        p10_mult_21_n410), .CO(p10_mult_21_n265), .S(p10_mult_21_n266) );
  FA_X1 p10_mult_21_U109 ( .A(p10_mult_21_n349), .B(p10_mult_21_n397), .CI(
        p10_mult_21_n373), .CO(p10_mult_21_n263), .S(p10_mult_21_n264) );
  FA_X1 p10_mult_21_U108 ( .A(p10_mult_21_n275), .B(p10_mult_21_n385), .CI(
        p10_mult_21_n273), .CO(p10_mult_21_n261), .S(p10_mult_21_n262) );
  FA_X1 p10_mult_21_U107 ( .A(p10_mult_21_n264), .B(p10_mult_21_n266), .CI(
        p10_mult_21_n271), .CO(p10_mult_21_n259), .S(p10_mult_21_n260) );
  FA_X1 p10_mult_21_U106 ( .A(p10_mult_21_n262), .B(p10_mult_21_n269), .CI(
        p10_mult_21_n260), .CO(p10_mult_21_n257), .S(p10_mult_21_n258) );
  HA_X1 p10_mult_21_U105 ( .A(p10_mult_21_n317), .B(p10_mult_21_n336), .CO(
        p10_mult_21_n255), .S(p10_mult_21_n256) );
  FA_X1 p10_mult_21_U104 ( .A(p10_mult_21_n409), .B(p10_mult_21_n372), .CI(
        p10_mult_21_n396), .CO(p10_mult_21_n253), .S(p10_mult_21_n254) );
  FA_X1 p10_mult_21_U103 ( .A(p10_mult_21_n348), .B(p10_mult_21_n384), .CI(
        p10_mult_21_n360), .CO(p10_mult_21_n251), .S(p10_mult_21_n252) );
  FA_X1 p10_mult_21_U102 ( .A(p10_mult_21_n265), .B(p10_mult_21_n256), .CI(
        p10_mult_21_n263), .CO(p10_mult_21_n249), .S(p10_mult_21_n250) );
  FA_X1 p10_mult_21_U101 ( .A(p10_mult_21_n254), .B(p10_mult_21_n252), .CI(
        p10_mult_21_n261), .CO(p10_mult_21_n247), .S(p10_mult_21_n248) );
  FA_X1 p10_mult_21_U100 ( .A(p10_mult_21_n259), .B(p10_mult_21_n250), .CI(
        p10_mult_21_n248), .CO(p10_mult_21_n245), .S(p10_mult_21_n246) );
  FA_X1 p10_mult_21_U97 ( .A(p10_mult_21_n395), .B(p10_mult_21_n359), .CI(
        p10_mult_21_n408), .CO(p10_mult_21_n241), .S(p10_mult_21_n242) );
  FA_X1 p10_mult_21_U96 ( .A(p10_mult_21_n335), .B(p10_mult_21_n371), .CI(
        p10_mult_21_n255), .CO(p10_mult_21_n239), .S(p10_mult_21_n240) );
  FA_X1 p10_mult_21_U95 ( .A(p10_mult_21_n253), .B(p10_mult_21_n244), .CI(
        p10_mult_21_n251), .CO(p10_mult_21_n237), .S(p10_mult_21_n238) );
  FA_X1 p10_mult_21_U94 ( .A(p10_mult_21_n240), .B(p10_mult_21_n242), .CI(
        p10_mult_21_n249), .CO(p10_mult_21_n235), .S(p10_mult_21_n236) );
  FA_X1 p10_mult_21_U93 ( .A(p10_mult_21_n247), .B(p10_mult_21_n238), .CI(
        p10_mult_21_n236), .CO(p10_mult_21_n233), .S(p10_mult_21_n234) );
  FA_X1 p10_mult_21_U91 ( .A(p10_mult_21_n382), .B(p10_mult_21_n346), .CI(
        p10_mult_21_n232), .CO(p10_mult_21_n229), .S(p10_mult_21_n230) );
  FA_X1 p10_mult_21_U90 ( .A(p10_mult_21_n334), .B(p10_mult_21_n370), .CI(
        p10_mult_21_n358), .CO(p10_mult_21_n227), .S(p10_mult_21_n228) );
  FA_X1 p10_mult_21_U89 ( .A(p10_mult_21_n241), .B(p10_mult_21_n243), .CI(
        p10_mult_21_n239), .CO(p10_mult_21_n225), .S(p10_mult_21_n226) );
  FA_X1 p10_mult_21_U88 ( .A(p10_mult_21_n230), .B(p10_mult_21_n228), .CI(
        p10_mult_21_n237), .CO(p10_mult_21_n223), .S(p10_mult_21_n224) );
  FA_X1 p10_mult_21_U87 ( .A(p10_mult_21_n235), .B(p10_mult_21_n226), .CI(
        p10_mult_21_n224), .CO(p10_mult_21_n221), .S(p10_mult_21_n222) );
  FA_X1 p10_mult_21_U86 ( .A(p10_mult_21_n231), .B(p10_mult_21_n333), .CI(
        p10_mult_21_n394), .CO(p10_mult_21_n219), .S(p10_mult_21_n220) );
  FA_X1 p10_mult_21_U85 ( .A(p10_mult_21_n345), .B(p10_mult_21_n381), .CI(
        p10_mult_21_n357), .CO(p10_mult_21_n217), .S(p10_mult_21_n218) );
  FA_X1 p10_mult_21_U84 ( .A(p10_mult_21_n229), .B(p10_mult_21_n369), .CI(
        p10_mult_21_n227), .CO(p10_mult_21_n215), .S(p10_mult_21_n216) );
  FA_X1 p10_mult_21_U83 ( .A(p10_mult_21_n220), .B(p10_mult_21_n218), .CI(
        p10_mult_21_n225), .CO(p10_mult_21_n213), .S(p10_mult_21_n214) );
  FA_X1 p10_mult_21_U82 ( .A(p10_mult_21_n223), .B(p10_mult_21_n216), .CI(
        p10_mult_21_n214), .CO(p10_mult_21_n211), .S(p10_mult_21_n212) );
  FA_X1 p10_mult_21_U80 ( .A(p10_mult_21_n368), .B(p10_mult_21_n344), .CI(
        p10_mult_21_n210), .CO(p10_mult_21_n207), .S(p10_mult_21_n208) );
  FA_X1 p10_mult_21_U79 ( .A(p10_mult_21_n332), .B(p10_mult_21_n356), .CI(
        p10_mult_21_n219), .CO(p10_mult_21_n205), .S(p10_mult_21_n206) );
  FA_X1 p10_mult_21_U78 ( .A(p10_mult_21_n208), .B(p10_mult_21_n217), .CI(
        p10_mult_21_n215), .CO(p10_mult_21_n203), .S(p10_mult_21_n204) );
  FA_X1 p10_mult_21_U77 ( .A(p10_mult_21_n213), .B(p10_mult_21_n206), .CI(
        p10_mult_21_n204), .CO(p10_mult_21_n201), .S(p10_mult_21_n202) );
  FA_X1 p10_mult_21_U76 ( .A(p10_mult_21_n209), .B(p10_mult_21_n331), .CI(
        p10_mult_21_n380), .CO(p10_mult_21_n199), .S(p10_mult_21_n200) );
  FA_X1 p10_mult_21_U75 ( .A(p10_mult_21_n355), .B(p10_mult_21_n343), .CI(
        p10_mult_21_n367), .CO(p10_mult_21_n197), .S(p10_mult_21_n198) );
  FA_X1 p10_mult_21_U74 ( .A(p10_mult_21_n198), .B(p10_mult_21_n207), .CI(
        p10_mult_21_n200), .CO(p10_mult_21_n195), .S(p10_mult_21_n196) );
  FA_X1 p10_mult_21_U73 ( .A(p10_mult_21_n203), .B(p10_mult_21_n205), .CI(
        p10_mult_21_n196), .CO(p10_mult_21_n193), .S(p10_mult_21_n194) );
  FA_X1 p10_mult_21_U71 ( .A(p10_mult_21_n330), .B(p10_mult_21_n342), .CI(
        p10_mult_21_n192), .CO(p10_mult_21_n189), .S(p10_mult_21_n190) );
  FA_X1 p10_mult_21_U70 ( .A(p10_mult_21_n199), .B(p10_mult_21_n354), .CI(
        p10_mult_21_n197), .CO(p10_mult_21_n187), .S(p10_mult_21_n188) );
  FA_X1 p10_mult_21_U69 ( .A(p10_mult_21_n188), .B(p10_mult_21_n190), .CI(
        p10_mult_21_n195), .CO(p10_mult_21_n185), .S(p10_mult_21_n186) );
  FA_X1 p10_mult_21_U68 ( .A(p10_mult_21_n191), .B(p10_mult_21_n329), .CI(
        p10_mult_21_n366), .CO(p10_mult_21_n183), .S(p10_mult_21_n184) );
  FA_X1 p10_mult_21_U67 ( .A(p10_mult_21_n341), .B(p10_mult_21_n353), .CI(
        p10_mult_21_n189), .CO(p10_mult_21_n181), .S(p10_mult_21_n182) );
  FA_X1 p10_mult_21_U66 ( .A(p10_mult_21_n187), .B(p10_mult_21_n184), .CI(
        p10_mult_21_n182), .CO(p10_mult_21_n179), .S(p10_mult_21_n180) );
  FA_X1 p10_mult_21_U64 ( .A(p10_mult_21_n328), .B(p10_mult_21_n340), .CI(
        p10_mult_21_n178), .CO(p10_mult_21_n175), .S(p10_mult_21_n176) );
  FA_X1 p10_mult_21_U63 ( .A(p10_mult_21_n176), .B(p10_mult_21_n183), .CI(
        p10_mult_21_n181), .CO(p10_mult_21_n173), .S(p10_mult_21_n174) );
  FA_X1 p10_mult_21_U62 ( .A(p10_mult_21_n327), .B(p10_mult_21_n177), .CI(
        p10_mult_21_n352), .CO(p10_mult_21_n171), .S(p10_mult_21_n172) );
  FA_X1 p10_mult_21_U61 ( .A(p10_mult_21_n175), .B(p10_mult_21_n339), .CI(
        p10_mult_21_n172), .CO(p10_mult_21_n169), .S(p10_mult_21_n170) );
  FA_X1 p10_mult_21_U59 ( .A(p10_mult_21_n168), .B(p10_mult_21_n326), .CI(
        p10_mult_21_n171), .CO(p10_mult_21_n165), .S(p10_mult_21_n166) );
  FA_X1 p10_mult_21_U58 ( .A(p10_mult_21_n325), .B(p10_mult_21_n167), .CI(
        p10_mult_21_n338), .CO(p10_mult_21_n163), .S(p10_mult_21_n164) );
  FA_X1 p10_mult_21_U44 ( .A(p10_mult_21_n246), .B(p10_mult_21_n257), .CI(
        p10_mult_21_n149), .CO(p10_mult_21_n148), .S(temp5[0]) );
  FA_X1 p10_mult_21_U43 ( .A(p10_mult_21_n234), .B(p10_mult_21_n245), .CI(
        p10_mult_21_n148), .CO(p10_mult_21_n147), .S(temp5[1]) );
  FA_X1 p10_mult_21_U42 ( .A(p10_mult_21_n222), .B(p10_mult_21_n233), .CI(
        p10_mult_21_n147), .CO(p10_mult_21_n146), .S(temp5[2]) );
  FA_X1 p10_mult_21_U41 ( .A(p10_mult_21_n212), .B(p10_mult_21_n221), .CI(
        p10_mult_21_n146), .CO(p10_mult_21_n145), .S(temp5[3]) );
  FA_X1 p10_mult_21_U40 ( .A(p10_mult_21_n202), .B(p10_mult_21_n211), .CI(
        p10_mult_21_n145), .CO(p10_mult_21_n144), .S(temp5[4]) );
  FA_X1 p10_mult_21_U39 ( .A(p10_mult_21_n194), .B(p10_mult_21_n201), .CI(
        p10_mult_21_n144), .CO(p10_mult_21_n143), .S(temp5[5]) );
  FA_X1 p10_mult_21_U38 ( .A(p10_mult_21_n186), .B(p10_mult_21_n193), .CI(
        p10_mult_21_n143), .CO(p10_mult_21_n142), .S(temp5[6]) );
  FA_X1 p10_mult_21_U37 ( .A(p10_mult_21_n180), .B(p10_mult_21_n185), .CI(
        p10_mult_21_n142), .CO(p10_mult_21_n141), .S(temp5[7]) );
  FA_X1 p10_mult_21_U30 ( .A(p10_mult_21_n174), .B(p10_mult_21_n179), .CI(
        p10_mult_21_n141), .CO(p10_mult_21_n140), .S(temp5[8]) );
  FA_X1 p10_mult_21_U20 ( .A(p10_mult_21_n170), .B(p10_mult_21_n173), .CI(
        p10_mult_21_n140), .CO(p10_mult_21_n139), .S(temp5[9]) );
  FA_X1 p10_mult_21_U10 ( .A(p10_mult_21_n166), .B(p10_mult_21_n169), .CI(
        p10_mult_21_n139), .CO(p10_mult_21_n138), .S(temp5[10]) );
  FA_X1 p10_mult_21_U9 ( .A(p10_mult_21_n165), .B(p10_mult_21_n164), .CI(
        p10_mult_21_n138), .CO(p10_mult_21_n137), .S(temp5[11]) );
  FA_X1 p10_mult_21_U8 ( .A(p10_mult_21_n163), .B(p10_mult_21_n162), .CI(
        p10_mult_21_n137), .CO(p10_mult_21_n136), .S(temp5[12]) );
  INV_X1 SUB1_U40 ( .A(reg7[0]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_1_) );
  INV_X1 SUB1_U39 ( .A(reg7[9]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_9_) );
  INV_X1 SUB1_U38 ( .A(reg7[8]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_8_) );
  INV_X1 SUB1_U37 ( .A(reg7[7]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_7_) );
  INV_X1 SUB1_U36 ( .A(reg7[6]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_6_) );
  INV_X1 SUB1_U35 ( .A(reg7[5]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_5_) );
  INV_X1 SUB1_U34 ( .A(reg7[4]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_4_) );
  INV_X1 SUB1_U33 ( .A(reg7[3]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_3_) );
  INV_X1 SUB1_U32 ( .A(reg7[2]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_2_) );
  INV_X1 SUB1_U31 ( .A(reg7[1]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_1_) );
  INV_X1 SUB1_U30 ( .A(reg7[13]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_13_) );
  INV_X1 SUB1_U29 ( .A(reg7[12]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_12_) );
  INV_X1 SUB1_U28 ( .A(reg7[11]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_11_) );
  INV_X1 SUB1_U27 ( .A(reg7[10]), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_10_) );
  XOR2_X1 SUB1_U26 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_1_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_1_), .Z(SUB1_N1) );
  AND2_X1 SUB1_U25 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_1_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_1_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_2_) );
  XOR2_X1 SUB1_U24 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_2_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_2_), .Z(SUB1_N2) );
  AND2_X1 SUB1_U23 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_2_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_2_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_3_) );
  XOR2_X1 SUB1_U22 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_3_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_3_), .Z(SUB1_N3) );
  AND2_X1 SUB1_U21 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_3_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_3_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_4_) );
  XOR2_X1 SUB1_U20 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_4_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_4_), .Z(SUB1_N4) );
  AND2_X1 SUB1_U19 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_4_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_4_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_5_) );
  XOR2_X1 SUB1_U18 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_5_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_5_), .Z(SUB1_N5) );
  AND2_X1 SUB1_U17 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_5_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_5_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_6_) );
  XOR2_X1 SUB1_U16 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_6_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_6_), .Z(SUB1_N6) );
  AND2_X1 SUB1_U15 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_6_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_6_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_7_) );
  XOR2_X1 SUB1_U14 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_7_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_7_), .Z(SUB1_N7) );
  AND2_X1 SUB1_U13 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_7_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_7_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_8_) );
  XOR2_X1 SUB1_U12 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_8_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_8_), .Z(SUB1_N8) );
  AND2_X1 SUB1_U11 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_8_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_8_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_9_) );
  XOR2_X1 SUB1_U10 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_9_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_9_), .Z(SUB1_N9) );
  AND2_X1 SUB1_U9 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_9_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_9_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_10_) );
  XOR2_X1 SUB1_U8 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_10_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_10_), .Z(SUB1_N10) );
  AND2_X1 SUB1_U7 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_10_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_10_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_11_) );
  XOR2_X1 SUB1_U6 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_11_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_11_), .Z(SUB1_N11) );
  AND2_X1 SUB1_U5 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_11_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_11_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_12_) );
  XOR2_X1 SUB1_U4 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_12_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_12_), .Z(SUB1_N12) );
  AND2_X1 SUB1_U3 ( .A1(SUB1_sub_1_root_sub_0_root_sub_21_2_carry_12_), .A2(
        SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_12_), .ZN(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_13_) );
  XOR2_X1 SUB1_U2 ( .A(SUB1_sub_1_root_sub_0_root_sub_21_2_B_not_13_), .B(
        SUB1_sub_1_root_sub_0_root_sub_21_2_carry_13_), .Z(SUB1_N13) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U16 ( .A(reg6[0]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U15 ( .A(reg6[10]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_10_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U14 ( .A(reg6[11]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U13 ( .A(reg6[12]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U12 ( .A(reg6[13]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_13_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U11 ( .A(reg6[1]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_1_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U10 ( .A(reg6[2]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_2_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U9 ( .A(reg6[3]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_3_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U8 ( .A(reg6[4]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_4_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U7 ( .A(reg6[5]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_5_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U6 ( .A(reg6[6]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_6_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U5 ( .A(reg6[7]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_7_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U4 ( .A(reg6[8]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_8_) );
  INV_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U3 ( .A(reg6[9]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_9_) );
  XNOR2_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2 ( .A(reg7[0]), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_), .ZN(fb[0]) );
  OR2_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U1 ( .A1(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_0_), .A2(reg7[0]), .ZN(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_1 ( .A(SUB1_N1), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_1_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_), .S(fb[1]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_2 ( .A(SUB1_N2), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_2_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_), .S(fb[2]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_3 ( .A(SUB1_N3), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_3_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_), .S(fb[3]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_4 ( .A(SUB1_N4), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_4_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_), .S(fb[4]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_5 ( .A(SUB1_N5), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_5_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_), .S(fb[5]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_6 ( .A(SUB1_N6), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_6_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_), .S(fb[6]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_7 ( .A(SUB1_N7), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_7_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_), .S(fb[7]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_8 ( .A(SUB1_N8), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_8_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_), .S(fb[8]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_9 ( .A(SUB1_N9), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_9_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_), .S(fb[9]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_10 ( .A(SUB1_N10), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_10_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_), .S(fb[10]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_11 ( .A(SUB1_N11), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_11_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_), .S(fb[11]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_12 ( .A(SUB1_N12), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_12_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_), .S(fb[12]) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_13 ( .A(SUB1_N13), .B(
        SUB1_sub_0_root_sub_0_root_sub_21_2_B_not_13_), .CI(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_), .S(fb[13]) );
  XOR2_X1 s6_add_21_U2 ( .A(mul2_reg[0]), .B(mul1_reg[0]), .Z(sig_ff1[0]) );
  AND2_X1 s6_add_21_U1 ( .A1(mul1_reg[0]), .A2(mul2_reg[0]), .ZN(
        s6_add_21_carry_1_) );
  FA_X1 s6_add_21_U1_1 ( .A(mul1_reg[1]), .B(mul2_reg[1]), .CI(
        s6_add_21_carry_1_), .CO(s6_add_21_carry_2_), .S(sig_ff1[1]) );
  FA_X1 s6_add_21_U1_2 ( .A(mul1_reg[2]), .B(mul2_reg[2]), .CI(
        s6_add_21_carry_2_), .CO(s6_add_21_carry_3_), .S(sig_ff1[2]) );
  FA_X1 s6_add_21_U1_3 ( .A(mul1_reg[3]), .B(mul2_reg[3]), .CI(
        s6_add_21_carry_3_), .CO(s6_add_21_carry_4_), .S(sig_ff1[3]) );
  FA_X1 s6_add_21_U1_4 ( .A(mul1_reg[4]), .B(mul2_reg[4]), .CI(
        s6_add_21_carry_4_), .CO(s6_add_21_carry_5_), .S(sig_ff1[4]) );
  FA_X1 s6_add_21_U1_5 ( .A(mul1_reg[5]), .B(mul2_reg[5]), .CI(
        s6_add_21_carry_5_), .CO(s6_add_21_carry_6_), .S(sig_ff1[5]) );
  FA_X1 s6_add_21_U1_6 ( .A(mul1_reg[6]), .B(mul2_reg[6]), .CI(
        s6_add_21_carry_6_), .CO(s6_add_21_carry_7_), .S(sig_ff1[6]) );
  FA_X1 s6_add_21_U1_7 ( .A(mul1_reg[7]), .B(mul2_reg[7]), .CI(
        s6_add_21_carry_7_), .CO(s6_add_21_carry_8_), .S(sig_ff1[7]) );
  FA_X1 s6_add_21_U1_8 ( .A(mul1_reg[8]), .B(mul2_reg[8]), .CI(
        s6_add_21_carry_8_), .CO(s6_add_21_carry_9_), .S(sig_ff1[8]) );
  FA_X1 s6_add_21_U1_9 ( .A(mul1_reg[9]), .B(mul2_reg[9]), .CI(
        s6_add_21_carry_9_), .CO(s6_add_21_carry_10_), .S(sig_ff1[9]) );
  FA_X1 s6_add_21_U1_10 ( .A(mul1_reg[10]), .B(mul2_reg[10]), .CI(
        s6_add_21_carry_10_), .CO(s6_add_21_carry_11_), .S(sig_ff1[10]) );
  FA_X1 s6_add_21_U1_11 ( .A(mul1_reg[11]), .B(mul2_reg[11]), .CI(
        s6_add_21_carry_11_), .CO(s6_add_21_carry_12_), .S(sig_ff1[11]) );
  FA_X1 s6_add_21_U1_12 ( .A(mul1_reg[12]), .B(mul2_reg[12]), .CI(
        s6_add_21_carry_12_), .CO(s6_add_21_carry_13_), .S(sig_ff1[12]) );
  FA_X1 s6_add_21_U1_13 ( .A(mul1_reg[13]), .B(mul2_reg[13]), .CI(
        s6_add_21_carry_13_), .S(sig_ff1[13]) );
  XOR2_X1 s7_add_21_U2 ( .A(mul4_reg[0]), .B(mul3_reg[0]), .Z(sig_ff2[0]) );
  AND2_X1 s7_add_21_U1 ( .A1(mul3_reg[0]), .A2(mul4_reg[0]), .ZN(
        s7_add_21_carry_1_) );
  FA_X1 s7_add_21_U1_1 ( .A(mul3_reg[1]), .B(mul4_reg[1]), .CI(
        s7_add_21_carry_1_), .CO(s7_add_21_carry_2_), .S(sig_ff2[1]) );
  FA_X1 s7_add_21_U1_2 ( .A(mul3_reg[2]), .B(mul4_reg[2]), .CI(
        s7_add_21_carry_2_), .CO(s7_add_21_carry_3_), .S(sig_ff2[2]) );
  FA_X1 s7_add_21_U1_3 ( .A(mul3_reg[3]), .B(mul4_reg[3]), .CI(
        s7_add_21_carry_3_), .CO(s7_add_21_carry_4_), .S(sig_ff2[3]) );
  FA_X1 s7_add_21_U1_4 ( .A(mul3_reg[4]), .B(mul4_reg[4]), .CI(
        s7_add_21_carry_4_), .CO(s7_add_21_carry_5_), .S(sig_ff2[4]) );
  FA_X1 s7_add_21_U1_5 ( .A(mul3_reg[5]), .B(mul4_reg[5]), .CI(
        s7_add_21_carry_5_), .CO(s7_add_21_carry_6_), .S(sig_ff2[5]) );
  FA_X1 s7_add_21_U1_6 ( .A(mul3_reg[6]), .B(mul4_reg[6]), .CI(
        s7_add_21_carry_6_), .CO(s7_add_21_carry_7_), .S(sig_ff2[6]) );
  FA_X1 s7_add_21_U1_7 ( .A(mul3_reg[7]), .B(mul4_reg[7]), .CI(
        s7_add_21_carry_7_), .CO(s7_add_21_carry_8_), .S(sig_ff2[7]) );
  FA_X1 s7_add_21_U1_8 ( .A(mul3_reg[8]), .B(mul4_reg[8]), .CI(
        s7_add_21_carry_8_), .CO(s7_add_21_carry_9_), .S(sig_ff2[8]) );
  FA_X1 s7_add_21_U1_9 ( .A(mul3_reg[9]), .B(mul4_reg[9]), .CI(
        s7_add_21_carry_9_), .CO(s7_add_21_carry_10_), .S(sig_ff2[9]) );
  FA_X1 s7_add_21_U1_10 ( .A(mul3_reg[10]), .B(mul4_reg[10]), .CI(
        s7_add_21_carry_10_), .CO(s7_add_21_carry_11_), .S(sig_ff2[10]) );
  FA_X1 s7_add_21_U1_11 ( .A(mul3_reg[11]), .B(mul4_reg[11]), .CI(
        s7_add_21_carry_11_), .CO(s7_add_21_carry_12_), .S(sig_ff2[11]) );
  FA_X1 s7_add_21_U1_12 ( .A(mul3_reg[12]), .B(mul4_reg[12]), .CI(
        s7_add_21_carry_12_), .CO(s7_add_21_carry_13_), .S(sig_ff2[12]) );
  FA_X1 s7_add_21_U1_13 ( .A(mul3_reg[13]), .B(mul4_reg[13]), .CI(
        s7_add_21_carry_13_), .S(sig_ff2[13]) );
  XOR2_X1 s8_add_21_U2 ( .A(sig_ff2[0]), .B(sig_ff1[0]), .Z(DOUT[0]) );
  AND2_X1 s8_add_21_U1 ( .A1(sig_ff1[0]), .A2(sig_ff2[0]), .ZN(
        s8_add_21_carry_1_) );
  FA_X1 s8_add_21_U1_1 ( .A(sig_ff1[1]), .B(sig_ff2[1]), .CI(
        s8_add_21_carry_1_), .CO(s8_add_21_carry_2_), .S(DOUT[1]) );
  FA_X1 s8_add_21_U1_2 ( .A(sig_ff1[2]), .B(sig_ff2[2]), .CI(
        s8_add_21_carry_2_), .CO(s8_add_21_carry_3_), .S(DOUT[2]) );
  FA_X1 s8_add_21_U1_3 ( .A(sig_ff1[3]), .B(sig_ff2[3]), .CI(
        s8_add_21_carry_3_), .CO(s8_add_21_carry_4_), .S(DOUT[3]) );
  FA_X1 s8_add_21_U1_4 ( .A(sig_ff1[4]), .B(sig_ff2[4]), .CI(
        s8_add_21_carry_4_), .CO(s8_add_21_carry_5_), .S(DOUT[4]) );
  FA_X1 s8_add_21_U1_5 ( .A(sig_ff1[5]), .B(sig_ff2[5]), .CI(
        s8_add_21_carry_5_), .CO(s8_add_21_carry_6_), .S(DOUT[5]) );
  FA_X1 s8_add_21_U1_6 ( .A(sig_ff1[6]), .B(sig_ff2[6]), .CI(
        s8_add_21_carry_6_), .CO(s8_add_21_carry_7_), .S(DOUT[6]) );
  FA_X1 s8_add_21_U1_7 ( .A(sig_ff1[7]), .B(sig_ff2[7]), .CI(
        s8_add_21_carry_7_), .CO(s8_add_21_carry_8_), .S(DOUT[7]) );
  FA_X1 s8_add_21_U1_8 ( .A(sig_ff1[8]), .B(sig_ff2[8]), .CI(
        s8_add_21_carry_8_), .CO(s8_add_21_carry_9_), .S(DOUT[8]) );
  FA_X1 s8_add_21_U1_9 ( .A(sig_ff1[9]), .B(sig_ff2[9]), .CI(
        s8_add_21_carry_9_), .CO(s8_add_21_carry_10_), .S(DOUT[9]) );
  FA_X1 s8_add_21_U1_10 ( .A(sig_ff1[10]), .B(sig_ff2[10]), .CI(
        s8_add_21_carry_10_), .CO(s8_add_21_carry_11_), .S(DOUT[10]) );
  FA_X1 s8_add_21_U1_11 ( .A(sig_ff1[11]), .B(sig_ff2[11]), .CI(
        s8_add_21_carry_11_), .CO(s8_add_21_carry_12_), .S(DOUT[11]) );
  FA_X1 s8_add_21_U1_12 ( .A(sig_ff1[12]), .B(sig_ff2[12]), .CI(
        s8_add_21_carry_12_), .CO(s8_add_21_carry_13_), .S(DOUT[12]) );
  FA_X1 s8_add_21_U1_13 ( .A(sig_ff1[13]), .B(sig_ff2[13]), .CI(
        s8_add_21_carry_13_), .S(DOUT[13]) );
  XOR2_X1 s9_add_21_U2 ( .A(xin[0]), .B(fb[0]), .Z(w[0]) );
  AND2_X1 s9_add_21_U1 ( .A1(fb[0]), .A2(xin[0]), .ZN(s9_add_21_carry_1_) );
  FA_X1 s9_add_21_U1_1 ( .A(fb[1]), .B(xin[1]), .CI(s9_add_21_carry_1_), .CO(
        s9_add_21_carry_2_), .S(w[1]) );
  FA_X1 s9_add_21_U1_2 ( .A(fb[2]), .B(xin[2]), .CI(s9_add_21_carry_2_), .CO(
        s9_add_21_carry_3_), .S(w[2]) );
  FA_X1 s9_add_21_U1_3 ( .A(fb[3]), .B(xin[3]), .CI(s9_add_21_carry_3_), .CO(
        s9_add_21_carry_4_), .S(w[3]) );
  FA_X1 s9_add_21_U1_4 ( .A(fb[4]), .B(xin[4]), .CI(s9_add_21_carry_4_), .CO(
        s9_add_21_carry_5_), .S(w[4]) );
  FA_X1 s9_add_21_U1_5 ( .A(fb[5]), .B(xin[5]), .CI(s9_add_21_carry_5_), .CO(
        s9_add_21_carry_6_), .S(w[5]) );
  FA_X1 s9_add_21_U1_6 ( .A(fb[6]), .B(xin[6]), .CI(s9_add_21_carry_6_), .CO(
        s9_add_21_carry_7_), .S(w[6]) );
  FA_X1 s9_add_21_U1_7 ( .A(fb[7]), .B(xin[7]), .CI(s9_add_21_carry_7_), .CO(
        s9_add_21_carry_8_), .S(w[7]) );
  FA_X1 s9_add_21_U1_8 ( .A(fb[8]), .B(xin[8]), .CI(s9_add_21_carry_8_), .CO(
        s9_add_21_carry_9_), .S(w[8]) );
  FA_X1 s9_add_21_U1_9 ( .A(fb[9]), .B(xin[9]), .CI(s9_add_21_carry_9_), .CO(
        s9_add_21_carry_10_), .S(w[9]) );
  FA_X1 s9_add_21_U1_10 ( .A(fb[10]), .B(xin[10]), .CI(s9_add_21_carry_10_), 
        .CO(s9_add_21_carry_11_), .S(w[10]) );
  FA_X1 s9_add_21_U1_11 ( .A(fb[11]), .B(xin[11]), .CI(s9_add_21_carry_11_), 
        .CO(s9_add_21_carry_12_), .S(w[11]) );
  FA_X1 s9_add_21_U1_12 ( .A(fb[12]), .B(xin[12]), .CI(s9_add_21_carry_12_), 
        .CO(s9_add_21_carry_13_), .S(w[12]) );
  FA_X1 s9_add_21_U1_13 ( .A(fb[13]), .B(xin[13]), .CI(s9_add_21_carry_13_), 
        .S(w[13]) );
  NAND2_X1 REG11_U34 ( .A1(w[13]), .A2(REG11_n43), .ZN(REG11_n76) );
  OAI21_X1 REG11_U33 ( .B1(REG11_n44), .B2(REG11_n75), .A(REG11_n76), .ZN(
        REG11_n48) );
  NAND2_X1 REG11_U32 ( .A1(w[6]), .A2(REG11_n43), .ZN(REG11_n83) );
  OAI21_X1 REG11_U31 ( .B1(REG11_n44), .B2(REG11_n68), .A(REG11_n83), .ZN(
        REG11_n55) );
  NAND2_X1 REG11_U30 ( .A1(w[5]), .A2(REG11_n43), .ZN(REG11_n84) );
  OAI21_X1 REG11_U29 ( .B1(REG11_n44), .B2(REG11_n67), .A(REG11_n84), .ZN(
        REG11_n56) );
  NAND2_X1 REG11_U28 ( .A1(w[4]), .A2(REG11_n43), .ZN(REG11_n85) );
  OAI21_X1 REG11_U27 ( .B1(REG11_n45), .B2(REG11_n66), .A(REG11_n85), .ZN(
        REG11_n57) );
  NAND2_X1 REG11_U26 ( .A1(w[3]), .A2(REG11_n43), .ZN(REG11_n86) );
  OAI21_X1 REG11_U25 ( .B1(REG11_n45), .B2(REG11_n65), .A(REG11_n86), .ZN(
        REG11_n58) );
  NAND2_X1 REG11_U24 ( .A1(w[2]), .A2(REG11_n43), .ZN(REG11_n87) );
  OAI21_X1 REG11_U23 ( .B1(REG11_n45), .B2(REG11_n64), .A(REG11_n87), .ZN(
        REG11_n59) );
  NAND2_X1 REG11_U22 ( .A1(w[1]), .A2(REG11_n43), .ZN(REG11_n88) );
  OAI21_X1 REG11_U21 ( .B1(REG11_n44), .B2(REG11_n63), .A(REG11_n88), .ZN(
        REG11_n60) );
  NAND2_X1 REG11_U20 ( .A1(w[8]), .A2(REG11_n44), .ZN(REG11_n81) );
  OAI21_X1 REG11_U19 ( .B1(REG11_n44), .B2(REG11_n70), .A(REG11_n81), .ZN(
        REG11_n53) );
  NAND2_X1 REG11_U18 ( .A1(w[12]), .A2(REG11_n43), .ZN(REG11_n77) );
  OAI21_X1 REG11_U17 ( .B1(REG11_n44), .B2(REG11_n74), .A(REG11_n77), .ZN(
        REG11_n49) );
  NAND2_X1 REG11_U16 ( .A1(w[11]), .A2(REG11_n43), .ZN(REG11_n78) );
  OAI21_X1 REG11_U15 ( .B1(REG11_n44), .B2(REG11_n73), .A(REG11_n78), .ZN(
        REG11_n50) );
  NAND2_X1 REG11_U14 ( .A1(w[10]), .A2(REG11_n44), .ZN(REG11_n79) );
  OAI21_X1 REG11_U13 ( .B1(REG11_n44), .B2(REG11_n72), .A(REG11_n79), .ZN(
        REG11_n51) );
  NAND2_X1 REG11_U12 ( .A1(w[9]), .A2(REG11_n43), .ZN(REG11_n80) );
  OAI21_X1 REG11_U11 ( .B1(REG11_n44), .B2(REG11_n71), .A(REG11_n80), .ZN(
        REG11_n52) );
  NAND2_X1 REG11_U10 ( .A1(w[7]), .A2(REG11_n43), .ZN(REG11_n82) );
  OAI21_X1 REG11_U9 ( .B1(REG11_n44), .B2(REG11_n69), .A(REG11_n82), .ZN(
        REG11_n54) );
  NAND2_X1 REG11_U8 ( .A1(w[0]), .A2(REG11_n43), .ZN(REG11_n89) );
  OAI21_X1 REG11_U7 ( .B1(REG11_n44), .B2(REG11_n62), .A(REG11_n89), .ZN(
        REG11_n61) );
  BUF_X1 REG11_U6 ( .A(n47), .Z(REG11_n47) );
  BUF_X1 REG11_U5 ( .A(n47), .Z(REG11_n46) );
  BUF_X1 REG11_U4 ( .A(VIN), .Z(REG11_n45) );
  BUF_X1 REG11_U3 ( .A(VIN), .Z(REG11_n43) );
  BUF_X1 REG11_U2 ( .A(VIN), .Z(REG11_n44) );
  DFFR_X1 REG11_q_reg_0_ ( .D(REG11_n61), .CK(CLK), .RN(REG11_n47), .Q(reg2[0]), .QN(REG11_n62) );
  DFFR_X1 REG11_q_reg_1_ ( .D(REG11_n60), .CK(CLK), .RN(REG11_n47), .Q(reg2[1]), .QN(REG11_n63) );
  DFFR_X1 REG11_q_reg_2_ ( .D(REG11_n59), .CK(CLK), .RN(REG11_n46), .Q(reg2[2]), .QN(REG11_n64) );
  DFFR_X1 REG11_q_reg_3_ ( .D(REG11_n58), .CK(CLK), .RN(REG11_n46), .Q(reg2[3]), .QN(REG11_n65) );
  DFFR_X1 REG11_q_reg_4_ ( .D(REG11_n57), .CK(CLK), .RN(REG11_n46), .Q(reg2[4]), .QN(REG11_n66) );
  DFFR_X1 REG11_q_reg_5_ ( .D(REG11_n56), .CK(CLK), .RN(REG11_n46), .Q(reg2[5]), .QN(REG11_n67) );
  DFFR_X1 REG11_q_reg_6_ ( .D(REG11_n55), .CK(CLK), .RN(REG11_n46), .Q(reg2[6]), .QN(REG11_n68) );
  DFFR_X1 REG11_q_reg_7_ ( .D(REG11_n54), .CK(CLK), .RN(REG11_n46), .Q(reg2[7]), .QN(REG11_n69) );
  DFFR_X1 REG11_q_reg_8_ ( .D(REG11_n53), .CK(CLK), .RN(REG11_n46), .Q(reg2[8]), .QN(REG11_n70) );
  DFFR_X1 REG11_q_reg_9_ ( .D(REG11_n52), .CK(CLK), .RN(REG11_n46), .Q(reg2[9]), .QN(REG11_n71) );
  DFFR_X1 REG11_q_reg_10_ ( .D(REG11_n51), .CK(CLK), .RN(REG11_n46), .Q(
        reg2[10]), .QN(REG11_n72) );
  DFFR_X1 REG11_q_reg_11_ ( .D(REG11_n50), .CK(CLK), .RN(REG11_n46), .Q(
        reg2[11]), .QN(REG11_n73) );
  DFFR_X1 REG11_q_reg_12_ ( .D(REG11_n49), .CK(CLK), .RN(REG11_n46), .Q(
        reg2[12]), .QN(REG11_n74) );
  DFFR_X1 REG11_q_reg_13_ ( .D(REG11_n48), .CK(CLK), .RN(REG11_n46), .Q(
        reg2[13]), .QN(REG11_n75) );
  NAND2_X1 REG21_U34 ( .A1(reg2[3]), .A2(REG21_n43), .ZN(REG21_n86) );
  OAI21_X1 REG21_U33 ( .B1(REG21_n45), .B2(REG21_n65), .A(REG21_n86), .ZN(
        REG21_n58) );
  NAND2_X1 REG21_U32 ( .A1(reg2[12]), .A2(REG21_n43), .ZN(REG21_n77) );
  OAI21_X1 REG21_U31 ( .B1(REG21_n44), .B2(REG21_n74), .A(REG21_n77), .ZN(
        REG21_n49) );
  NAND2_X1 REG21_U30 ( .A1(reg2[6]), .A2(REG21_n43), .ZN(REG21_n83) );
  OAI21_X1 REG21_U29 ( .B1(REG21_n44), .B2(REG21_n68), .A(REG21_n83), .ZN(
        REG21_n55) );
  NAND2_X1 REG21_U28 ( .A1(reg2[4]), .A2(REG21_n43), .ZN(REG21_n85) );
  OAI21_X1 REG21_U27 ( .B1(REG21_n45), .B2(REG21_n66), .A(REG21_n85), .ZN(
        REG21_n57) );
  NAND2_X1 REG21_U26 ( .A1(reg2[2]), .A2(REG21_n43), .ZN(REG21_n87) );
  OAI21_X1 REG21_U25 ( .B1(REG21_n45), .B2(REG21_n64), .A(REG21_n87), .ZN(
        REG21_n59) );
  NAND2_X1 REG21_U24 ( .A1(reg2[0]), .A2(REG21_n43), .ZN(REG21_n89) );
  OAI21_X1 REG21_U23 ( .B1(REG21_n44), .B2(REG21_n62), .A(REG21_n89), .ZN(
        REG21_n61) );
  NAND2_X1 REG21_U22 ( .A1(reg2[13]), .A2(REG21_n43), .ZN(REG21_n76) );
  OAI21_X1 REG21_U21 ( .B1(REG21_n44), .B2(REG21_n75), .A(REG21_n76), .ZN(
        REG21_n48) );
  NAND2_X1 REG21_U20 ( .A1(reg2[10]), .A2(REG21_n44), .ZN(REG21_n79) );
  OAI21_X1 REG21_U19 ( .B1(REG21_n44), .B2(REG21_n72), .A(REG21_n79), .ZN(
        REG21_n51) );
  NAND2_X1 REG21_U18 ( .A1(reg2[8]), .A2(REG21_n44), .ZN(REG21_n81) );
  OAI21_X1 REG21_U17 ( .B1(REG21_n44), .B2(REG21_n70), .A(REG21_n81), .ZN(
        REG21_n53) );
  NAND2_X1 REG21_U16 ( .A1(reg2[1]), .A2(REG21_n43), .ZN(REG21_n88) );
  OAI21_X1 REG21_U15 ( .B1(REG21_n44), .B2(REG21_n63), .A(REG21_n88), .ZN(
        REG21_n60) );
  NAND2_X1 REG21_U14 ( .A1(reg2[11]), .A2(REG21_n43), .ZN(REG21_n78) );
  OAI21_X1 REG21_U13 ( .B1(REG21_n44), .B2(REG21_n73), .A(REG21_n78), .ZN(
        REG21_n50) );
  NAND2_X1 REG21_U12 ( .A1(reg2[9]), .A2(REG21_n43), .ZN(REG21_n80) );
  OAI21_X1 REG21_U11 ( .B1(REG21_n44), .B2(REG21_n71), .A(REG21_n80), .ZN(
        REG21_n52) );
  NAND2_X1 REG21_U10 ( .A1(reg2[7]), .A2(REG21_n43), .ZN(REG21_n82) );
  OAI21_X1 REG21_U9 ( .B1(REG21_n44), .B2(REG21_n69), .A(REG21_n82), .ZN(
        REG21_n54) );
  NAND2_X1 REG21_U8 ( .A1(reg2[5]), .A2(REG21_n43), .ZN(REG21_n84) );
  OAI21_X1 REG21_U7 ( .B1(REG21_n44), .B2(REG21_n67), .A(REG21_n84), .ZN(
        REG21_n56) );
  BUF_X1 REG21_U6 ( .A(n47), .Z(REG21_n47) );
  BUF_X1 REG21_U5 ( .A(n47), .Z(REG21_n46) );
  BUF_X1 REG21_U4 ( .A(VIN), .Z(REG21_n45) );
  BUF_X1 REG21_U3 ( .A(VIN), .Z(REG21_n43) );
  BUF_X1 REG21_U2 ( .A(VIN), .Z(REG21_n44) );
  DFFR_X1 REG21_q_reg_0_ ( .D(REG21_n61), .CK(CLK), .RN(REG21_n47), .Q(reg3[0]), .QN(REG21_n62) );
  DFFR_X1 REG21_q_reg_1_ ( .D(REG21_n60), .CK(CLK), .RN(REG21_n47), .Q(reg3[1]), .QN(REG21_n63) );
  DFFR_X1 REG21_q_reg_2_ ( .D(REG21_n59), .CK(CLK), .RN(REG21_n46), .Q(reg3[2]), .QN(REG21_n64) );
  DFFR_X1 REG21_q_reg_3_ ( .D(REG21_n58), .CK(CLK), .RN(REG21_n46), .Q(reg3[3]), .QN(REG21_n65) );
  DFFR_X1 REG21_q_reg_4_ ( .D(REG21_n57), .CK(CLK), .RN(REG21_n46), .Q(reg3[4]), .QN(REG21_n66) );
  DFFR_X1 REG21_q_reg_5_ ( .D(REG21_n56), .CK(CLK), .RN(REG21_n46), .Q(reg3[5]), .QN(REG21_n67) );
  DFFR_X1 REG21_q_reg_6_ ( .D(REG21_n55), .CK(CLK), .RN(REG21_n46), .Q(reg3[6]), .QN(REG21_n68) );
  DFFR_X1 REG21_q_reg_7_ ( .D(REG21_n54), .CK(CLK), .RN(REG21_n46), .Q(reg3[7]), .QN(REG21_n69) );
  DFFR_X1 REG21_q_reg_8_ ( .D(REG21_n53), .CK(CLK), .RN(REG21_n46), .Q(reg3[8]), .QN(REG21_n70) );
  DFFR_X1 REG21_q_reg_9_ ( .D(REG21_n52), .CK(CLK), .RN(REG21_n46), .Q(reg3[9]), .QN(REG21_n71) );
  DFFR_X1 REG21_q_reg_10_ ( .D(REG21_n51), .CK(CLK), .RN(REG21_n46), .Q(
        reg3[10]), .QN(REG21_n72) );
  DFFR_X1 REG21_q_reg_11_ ( .D(REG21_n50), .CK(CLK), .RN(REG21_n46), .Q(
        reg3[11]), .QN(REG21_n73) );
  DFFR_X1 REG21_q_reg_12_ ( .D(REG21_n49), .CK(CLK), .RN(REG21_n46), .Q(
        reg3[12]), .QN(REG21_n74) );
  DFFR_X1 REG21_q_reg_13_ ( .D(REG21_n48), .CK(CLK), .RN(REG21_n46), .Q(
        reg3[13]), .QN(REG21_n75) );
  NAND2_X1 REG31_U34 ( .A1(reg2[3]), .A2(REG31_n43), .ZN(REG31_n86) );
  OAI21_X1 REG31_U33 ( .B1(REG31_n45), .B2(REG31_n65), .A(REG31_n86), .ZN(
        REG31_n58) );
  NAND2_X1 REG31_U32 ( .A1(reg2[12]), .A2(REG31_n43), .ZN(REG31_n77) );
  OAI21_X1 REG31_U31 ( .B1(REG31_n44), .B2(REG31_n74), .A(REG31_n77), .ZN(
        REG31_n49) );
  NAND2_X1 REG31_U30 ( .A1(reg2[6]), .A2(REG31_n43), .ZN(REG31_n83) );
  OAI21_X1 REG31_U29 ( .B1(REG31_n44), .B2(REG31_n68), .A(REG31_n83), .ZN(
        REG31_n55) );
  NAND2_X1 REG31_U28 ( .A1(reg2[4]), .A2(REG31_n43), .ZN(REG31_n85) );
  OAI21_X1 REG31_U27 ( .B1(REG31_n45), .B2(REG31_n66), .A(REG31_n85), .ZN(
        REG31_n57) );
  NAND2_X1 REG31_U26 ( .A1(reg2[2]), .A2(REG31_n43), .ZN(REG31_n87) );
  OAI21_X1 REG31_U25 ( .B1(REG31_n45), .B2(REG31_n64), .A(REG31_n87), .ZN(
        REG31_n59) );
  NAND2_X1 REG31_U24 ( .A1(reg2[0]), .A2(REG31_n43), .ZN(REG31_n89) );
  OAI21_X1 REG31_U23 ( .B1(REG31_n44), .B2(REG31_n62), .A(REG31_n89), .ZN(
        REG31_n61) );
  NAND2_X1 REG31_U22 ( .A1(reg2[13]), .A2(REG31_n43), .ZN(REG31_n76) );
  OAI21_X1 REG31_U21 ( .B1(REG31_n44), .B2(REG31_n75), .A(REG31_n76), .ZN(
        REG31_n48) );
  NAND2_X1 REG31_U20 ( .A1(reg2[10]), .A2(REG31_n44), .ZN(REG31_n79) );
  OAI21_X1 REG31_U19 ( .B1(REG31_n44), .B2(REG31_n72), .A(REG31_n79), .ZN(
        REG31_n51) );
  NAND2_X1 REG31_U18 ( .A1(reg2[8]), .A2(REG31_n44), .ZN(REG31_n81) );
  OAI21_X1 REG31_U17 ( .B1(REG31_n44), .B2(REG31_n70), .A(REG31_n81), .ZN(
        REG31_n53) );
  NAND2_X1 REG31_U16 ( .A1(reg2[1]), .A2(REG31_n43), .ZN(REG31_n88) );
  OAI21_X1 REG31_U15 ( .B1(REG31_n44), .B2(REG31_n63), .A(REG31_n88), .ZN(
        REG31_n60) );
  NAND2_X1 REG31_U14 ( .A1(reg2[11]), .A2(REG31_n43), .ZN(REG31_n78) );
  OAI21_X1 REG31_U13 ( .B1(REG31_n44), .B2(REG31_n73), .A(REG31_n78), .ZN(
        REG31_n50) );
  NAND2_X1 REG31_U12 ( .A1(reg2[9]), .A2(REG31_n43), .ZN(REG31_n80) );
  OAI21_X1 REG31_U11 ( .B1(REG31_n44), .B2(REG31_n71), .A(REG31_n80), .ZN(
        REG31_n52) );
  NAND2_X1 REG31_U10 ( .A1(reg2[7]), .A2(REG31_n43), .ZN(REG31_n82) );
  OAI21_X1 REG31_U9 ( .B1(REG31_n44), .B2(REG31_n69), .A(REG31_n82), .ZN(
        REG31_n54) );
  NAND2_X1 REG31_U8 ( .A1(reg2[5]), .A2(REG31_n43), .ZN(REG31_n84) );
  OAI21_X1 REG31_U7 ( .B1(REG31_n44), .B2(REG31_n67), .A(REG31_n84), .ZN(
        REG31_n56) );
  BUF_X1 REG31_U6 ( .A(n47), .Z(REG31_n47) );
  BUF_X1 REG31_U5 ( .A(n47), .Z(REG31_n46) );
  BUF_X1 REG31_U4 ( .A(VIN), .Z(REG31_n45) );
  BUF_X1 REG31_U3 ( .A(VIN), .Z(REG31_n43) );
  BUF_X1 REG31_U2 ( .A(VIN), .Z(REG31_n44) );
  DFFR_X1 REG31_q_reg_0_ ( .D(REG31_n61), .CK(CLK), .RN(REG31_n47), .Q(reg4[0]), .QN(REG31_n62) );
  DFFR_X1 REG31_q_reg_1_ ( .D(REG31_n60), .CK(CLK), .RN(REG31_n47), .Q(reg4[1]), .QN(REG31_n63) );
  DFFR_X1 REG31_q_reg_2_ ( .D(REG31_n59), .CK(CLK), .RN(REG31_n46), .Q(reg4[2]), .QN(REG31_n64) );
  DFFR_X1 REG31_q_reg_3_ ( .D(REG31_n58), .CK(CLK), .RN(REG31_n46), .Q(reg4[3]), .QN(REG31_n65) );
  DFFR_X1 REG31_q_reg_4_ ( .D(REG31_n57), .CK(CLK), .RN(REG31_n46), .Q(reg4[4]), .QN(REG31_n66) );
  DFFR_X1 REG31_q_reg_5_ ( .D(REG31_n56), .CK(CLK), .RN(REG31_n46), .Q(reg4[5]), .QN(REG31_n67) );
  DFFR_X1 REG31_q_reg_6_ ( .D(REG31_n55), .CK(CLK), .RN(REG31_n46), .Q(reg4[6]), .QN(REG31_n68) );
  DFFR_X1 REG31_q_reg_7_ ( .D(REG31_n54), .CK(CLK), .RN(REG31_n46), .Q(reg4[7]), .QN(REG31_n69) );
  DFFR_X1 REG31_q_reg_8_ ( .D(REG31_n53), .CK(CLK), .RN(REG31_n46), .Q(reg4[8]), .QN(REG31_n70) );
  DFFR_X1 REG31_q_reg_9_ ( .D(REG31_n52), .CK(CLK), .RN(REG31_n46), .Q(reg4[9]), .QN(REG31_n71) );
  DFFR_X1 REG31_q_reg_10_ ( .D(REG31_n51), .CK(CLK), .RN(REG31_n46), .Q(
        reg4[10]), .QN(REG31_n72) );
  DFFR_X1 REG31_q_reg_11_ ( .D(REG31_n50), .CK(CLK), .RN(REG31_n46), .Q(
        reg4[11]), .QN(REG31_n73) );
  DFFR_X1 REG31_q_reg_12_ ( .D(REG31_n49), .CK(CLK), .RN(REG31_n46), .Q(
        reg4[12]), .QN(REG31_n74) );
  DFFR_X1 REG31_q_reg_13_ ( .D(REG31_n48), .CK(CLK), .RN(REG31_n46), .Q(
        reg4[13]), .QN(REG31_n75) );
  NAND2_X1 REG41_U34 ( .A1(reg4[4]), .A2(REG41_n43), .ZN(REG41_n85) );
  OAI21_X1 REG41_U33 ( .B1(REG41_n45), .B2(REG41_n66), .A(REG41_n85), .ZN(
        REG41_n57) );
  NAND2_X1 REG41_U32 ( .A1(reg4[2]), .A2(REG41_n43), .ZN(REG41_n87) );
  OAI21_X1 REG41_U31 ( .B1(REG41_n45), .B2(REG41_n64), .A(REG41_n87), .ZN(
        REG41_n59) );
  NAND2_X1 REG41_U30 ( .A1(reg4[0]), .A2(REG41_n43), .ZN(REG41_n89) );
  OAI21_X1 REG41_U29 ( .B1(REG41_n44), .B2(REG41_n62), .A(REG41_n89), .ZN(
        REG41_n61) );
  NAND2_X1 REG41_U28 ( .A1(reg4[13]), .A2(REG41_n43), .ZN(REG41_n76) );
  OAI21_X1 REG41_U27 ( .B1(REG41_n44), .B2(REG41_n75), .A(REG41_n76), .ZN(
        REG41_n48) );
  NAND2_X1 REG41_U26 ( .A1(reg4[12]), .A2(REG41_n43), .ZN(REG41_n77) );
  OAI21_X1 REG41_U25 ( .B1(REG41_n44), .B2(REG41_n74), .A(REG41_n77), .ZN(
        REG41_n49) );
  NAND2_X1 REG41_U24 ( .A1(reg4[10]), .A2(REG41_n44), .ZN(REG41_n79) );
  OAI21_X1 REG41_U23 ( .B1(REG41_n44), .B2(REG41_n72), .A(REG41_n79), .ZN(
        REG41_n51) );
  NAND2_X1 REG41_U22 ( .A1(reg4[8]), .A2(REG41_n44), .ZN(REG41_n81) );
  OAI21_X1 REG41_U21 ( .B1(REG41_n44), .B2(REG41_n70), .A(REG41_n81), .ZN(
        REG41_n53) );
  NAND2_X1 REG41_U20 ( .A1(reg4[6]), .A2(REG41_n43), .ZN(REG41_n83) );
  OAI21_X1 REG41_U19 ( .B1(REG41_n44), .B2(REG41_n68), .A(REG41_n83), .ZN(
        REG41_n55) );
  NAND2_X1 REG41_U18 ( .A1(reg4[1]), .A2(REG41_n43), .ZN(REG41_n88) );
  OAI21_X1 REG41_U17 ( .B1(REG41_n44), .B2(REG41_n63), .A(REG41_n88), .ZN(
        REG41_n60) );
  NAND2_X1 REG41_U16 ( .A1(reg4[11]), .A2(REG41_n43), .ZN(REG41_n78) );
  OAI21_X1 REG41_U15 ( .B1(REG41_n44), .B2(REG41_n73), .A(REG41_n78), .ZN(
        REG41_n50) );
  NAND2_X1 REG41_U14 ( .A1(reg4[9]), .A2(REG41_n43), .ZN(REG41_n80) );
  OAI21_X1 REG41_U13 ( .B1(REG41_n44), .B2(REG41_n71), .A(REG41_n80), .ZN(
        REG41_n52) );
  NAND2_X1 REG41_U12 ( .A1(reg4[7]), .A2(REG41_n43), .ZN(REG41_n82) );
  OAI21_X1 REG41_U11 ( .B1(REG41_n44), .B2(REG41_n69), .A(REG41_n82), .ZN(
        REG41_n54) );
  NAND2_X1 REG41_U10 ( .A1(reg4[5]), .A2(REG41_n43), .ZN(REG41_n84) );
  OAI21_X1 REG41_U9 ( .B1(REG41_n44), .B2(REG41_n67), .A(REG41_n84), .ZN(
        REG41_n56) );
  NAND2_X1 REG41_U8 ( .A1(reg4[3]), .A2(REG41_n43), .ZN(REG41_n86) );
  OAI21_X1 REG41_U7 ( .B1(REG41_n45), .B2(REG41_n65), .A(REG41_n86), .ZN(
        REG41_n58) );
  BUF_X1 REG41_U6 ( .A(n47), .Z(REG41_n47) );
  BUF_X1 REG41_U5 ( .A(n47), .Z(REG41_n46) );
  BUF_X1 REG41_U4 ( .A(VIN), .Z(REG41_n45) );
  BUF_X1 REG41_U3 ( .A(VIN), .Z(REG41_n43) );
  BUF_X1 REG41_U2 ( .A(VIN), .Z(REG41_n44) );
  DFFR_X1 REG41_q_reg_0_ ( .D(REG41_n61), .CK(CLK), .RN(REG41_n47), .Q(reg5[0]), .QN(REG41_n62) );
  DFFR_X1 REG41_q_reg_1_ ( .D(REG41_n60), .CK(CLK), .RN(REG41_n47), .Q(reg5[1]), .QN(REG41_n63) );
  DFFR_X1 REG41_q_reg_2_ ( .D(REG41_n59), .CK(CLK), .RN(REG41_n46), .Q(reg5[2]), .QN(REG41_n64) );
  DFFR_X1 REG41_q_reg_3_ ( .D(REG41_n58), .CK(CLK), .RN(REG41_n46), .Q(reg5[3]), .QN(REG41_n65) );
  DFFR_X1 REG41_q_reg_4_ ( .D(REG41_n57), .CK(CLK), .RN(REG41_n46), .Q(reg5[4]), .QN(REG41_n66) );
  DFFR_X1 REG41_q_reg_5_ ( .D(REG41_n56), .CK(CLK), .RN(REG41_n46), .Q(reg5[5]), .QN(REG41_n67) );
  DFFR_X1 REG41_q_reg_6_ ( .D(REG41_n55), .CK(CLK), .RN(REG41_n46), .Q(reg5[6]), .QN(REG41_n68) );
  DFFR_X1 REG41_q_reg_7_ ( .D(REG41_n54), .CK(CLK), .RN(REG41_n46), .Q(reg5[7]), .QN(REG41_n69) );
  DFFR_X1 REG41_q_reg_8_ ( .D(REG41_n53), .CK(CLK), .RN(REG41_n46), .Q(reg5[8]), .QN(REG41_n70) );
  DFFR_X1 REG41_q_reg_9_ ( .D(REG41_n52), .CK(CLK), .RN(REG41_n46), .Q(reg5[9]), .QN(REG41_n71) );
  DFFR_X1 REG41_q_reg_10_ ( .D(REG41_n51), .CK(CLK), .RN(REG41_n46), .Q(
        reg5[10]), .QN(REG41_n72) );
  DFFR_X1 REG41_q_reg_11_ ( .D(REG41_n50), .CK(CLK), .RN(REG41_n46), .Q(
        reg5[11]), .QN(REG41_n73) );
  DFFR_X1 REG41_q_reg_12_ ( .D(REG41_n49), .CK(CLK), .RN(REG41_n46), .Q(
        reg5[12]), .QN(REG41_n74) );
  DFFR_X1 REG41_q_reg_13_ ( .D(REG41_n48), .CK(CLK), .RN(REG41_n46), .Q(
        reg5[13]), .QN(REG41_n75) );
  NAND2_X1 REG51_U34 ( .A1(temp5[3]), .A2(REG51_n43), .ZN(REG51_n86) );
  OAI21_X1 REG51_U33 ( .B1(REG51_n45), .B2(REG51_n65), .A(REG51_n86), .ZN(
        REG51_n58) );
  NAND2_X1 REG51_U32 ( .A1(temp5[2]), .A2(REG51_n43), .ZN(REG51_n87) );
  OAI21_X1 REG51_U31 ( .B1(REG51_n45), .B2(REG51_n64), .A(REG51_n87), .ZN(
        REG51_n59) );
  NAND2_X1 REG51_U30 ( .A1(temp5[7]), .A2(REG51_n43), .ZN(REG51_n82) );
  OAI21_X1 REG51_U29 ( .B1(REG51_n44), .B2(REG51_n69), .A(REG51_n82), .ZN(
        REG51_n54) );
  NAND2_X1 REG51_U28 ( .A1(temp5[4]), .A2(REG51_n43), .ZN(REG51_n85) );
  OAI21_X1 REG51_U27 ( .B1(REG51_n45), .B2(REG51_n66), .A(REG51_n85), .ZN(
        REG51_n57) );
  NAND2_X1 REG51_U26 ( .A1(temp5[8]), .A2(REG51_n44), .ZN(REG51_n81) );
  OAI21_X1 REG51_U25 ( .B1(REG51_n44), .B2(REG51_n70), .A(REG51_n81), .ZN(
        REG51_n53) );
  NAND2_X1 REG51_U24 ( .A1(temp5[9]), .A2(REG51_n43), .ZN(REG51_n80) );
  OAI21_X1 REG51_U23 ( .B1(REG51_n44), .B2(REG51_n71), .A(REG51_n80), .ZN(
        REG51_n52) );
  NAND2_X1 REG51_U22 ( .A1(temp5[6]), .A2(REG51_n43), .ZN(REG51_n83) );
  OAI21_X1 REG51_U21 ( .B1(REG51_n44), .B2(REG51_n68), .A(REG51_n83), .ZN(
        REG51_n55) );
  NAND2_X1 REG51_U20 ( .A1(temp5[5]), .A2(REG51_n43), .ZN(REG51_n84) );
  OAI21_X1 REG51_U19 ( .B1(REG51_n44), .B2(REG51_n67), .A(REG51_n84), .ZN(
        REG51_n56) );
  NAND2_X1 REG51_U18 ( .A1(temp5[1]), .A2(REG51_n43), .ZN(REG51_n88) );
  OAI21_X1 REG51_U17 ( .B1(REG51_n44), .B2(REG51_n63), .A(REG51_n88), .ZN(
        REG51_n60) );
  NAND2_X1 REG51_U16 ( .A1(temp5[0]), .A2(REG51_n43), .ZN(REG51_n89) );
  OAI21_X1 REG51_U15 ( .B1(REG51_n44), .B2(REG51_n62), .A(REG51_n89), .ZN(
        REG51_n61) );
  NAND2_X1 REG51_U14 ( .A1(temp5[13]), .A2(REG51_n43), .ZN(REG51_n76) );
  OAI21_X1 REG51_U13 ( .B1(REG51_n44), .B2(REG51_n75), .A(REG51_n76), .ZN(
        REG51_n48) );
  NAND2_X1 REG51_U12 ( .A1(temp5[12]), .A2(REG51_n43), .ZN(REG51_n77) );
  OAI21_X1 REG51_U11 ( .B1(REG51_n44), .B2(REG51_n74), .A(REG51_n77), .ZN(
        REG51_n49) );
  NAND2_X1 REG51_U10 ( .A1(temp5[11]), .A2(REG51_n43), .ZN(REG51_n78) );
  OAI21_X1 REG51_U9 ( .B1(REG51_n44), .B2(REG51_n73), .A(REG51_n78), .ZN(
        REG51_n50) );
  NAND2_X1 REG51_U8 ( .A1(temp5[10]), .A2(REG51_n44), .ZN(REG51_n79) );
  OAI21_X1 REG51_U7 ( .B1(REG51_n44), .B2(REG51_n72), .A(REG51_n79), .ZN(
        REG51_n51) );
  BUF_X1 REG51_U6 ( .A(n47), .Z(REG51_n47) );
  BUF_X1 REG51_U5 ( .A(n47), .Z(REG51_n46) );
  BUF_X1 REG51_U4 ( .A(VIN), .Z(REG51_n45) );
  BUF_X1 REG51_U3 ( .A(VIN), .Z(REG51_n43) );
  BUF_X1 REG51_U2 ( .A(VIN), .Z(REG51_n44) );
  DFFR_X1 REG51_q_reg_0_ ( .D(REG51_n61), .CK(CLK), .RN(REG51_n47), .Q(reg6[0]), .QN(REG51_n62) );
  DFFR_X1 REG51_q_reg_1_ ( .D(REG51_n60), .CK(CLK), .RN(REG51_n47), .Q(reg6[1]), .QN(REG51_n63) );
  DFFR_X1 REG51_q_reg_2_ ( .D(REG51_n59), .CK(CLK), .RN(REG51_n46), .Q(reg6[2]), .QN(REG51_n64) );
  DFFR_X1 REG51_q_reg_3_ ( .D(REG51_n58), .CK(CLK), .RN(REG51_n46), .Q(reg6[3]), .QN(REG51_n65) );
  DFFR_X1 REG51_q_reg_4_ ( .D(REG51_n57), .CK(CLK), .RN(REG51_n46), .Q(reg6[4]), .QN(REG51_n66) );
  DFFR_X1 REG51_q_reg_5_ ( .D(REG51_n56), .CK(CLK), .RN(REG51_n46), .Q(reg6[5]), .QN(REG51_n67) );
  DFFR_X1 REG51_q_reg_6_ ( .D(REG51_n55), .CK(CLK), .RN(REG51_n46), .Q(reg6[6]), .QN(REG51_n68) );
  DFFR_X1 REG51_q_reg_7_ ( .D(REG51_n54), .CK(CLK), .RN(REG51_n46), .Q(reg6[7]), .QN(REG51_n69) );
  DFFR_X1 REG51_q_reg_8_ ( .D(REG51_n53), .CK(CLK), .RN(REG51_n46), .Q(reg6[8]), .QN(REG51_n70) );
  DFFR_X1 REG51_q_reg_9_ ( .D(REG51_n52), .CK(CLK), .RN(REG51_n46), .Q(reg6[9]), .QN(REG51_n71) );
  DFFR_X1 REG51_q_reg_10_ ( .D(REG51_n51), .CK(CLK), .RN(REG51_n46), .Q(
        reg6[10]), .QN(REG51_n72) );
  DFFR_X1 REG51_q_reg_11_ ( .D(REG51_n50), .CK(CLK), .RN(REG51_n46), .Q(
        reg6[11]), .QN(REG51_n73) );
  DFFR_X1 REG51_q_reg_12_ ( .D(REG51_n49), .CK(CLK), .RN(REG51_n46), .Q(
        reg6[12]), .QN(REG51_n74) );
  DFFR_X1 REG51_q_reg_13_ ( .D(REG51_n48), .CK(CLK), .RN(REG51_n46), .Q(
        reg6[13]), .QN(REG51_n75) );
  NAND2_X1 REG61_U34 ( .A1(temp6[4]), .A2(REG61_n43), .ZN(REG61_n85) );
  OAI21_X1 REG61_U33 ( .B1(REG61_n45), .B2(REG61_n66), .A(REG61_n85), .ZN(
        REG61_n57) );
  NAND2_X1 REG61_U32 ( .A1(temp6[2]), .A2(REG61_n43), .ZN(REG61_n87) );
  OAI21_X1 REG61_U31 ( .B1(REG61_n45), .B2(REG61_n64), .A(REG61_n87), .ZN(
        REG61_n59) );
  NAND2_X1 REG61_U30 ( .A1(temp6[3]), .A2(REG61_n43), .ZN(REG61_n86) );
  OAI21_X1 REG61_U29 ( .B1(REG61_n45), .B2(REG61_n65), .A(REG61_n86), .ZN(
        REG61_n58) );
  NAND2_X1 REG61_U28 ( .A1(temp6[8]), .A2(REG61_n44), .ZN(REG61_n81) );
  OAI21_X1 REG61_U27 ( .B1(REG61_n44), .B2(REG61_n70), .A(REG61_n81), .ZN(
        REG61_n53) );
  NAND2_X1 REG61_U26 ( .A1(temp6[9]), .A2(REG61_n43), .ZN(REG61_n80) );
  OAI21_X1 REG61_U25 ( .B1(REG61_n44), .B2(REG61_n71), .A(REG61_n80), .ZN(
        REG61_n52) );
  NAND2_X1 REG61_U24 ( .A1(temp6[7]), .A2(REG61_n43), .ZN(REG61_n82) );
  OAI21_X1 REG61_U23 ( .B1(REG61_n44), .B2(REG61_n69), .A(REG61_n82), .ZN(
        REG61_n54) );
  NAND2_X1 REG61_U22 ( .A1(temp6[6]), .A2(REG61_n43), .ZN(REG61_n83) );
  OAI21_X1 REG61_U21 ( .B1(REG61_n44), .B2(REG61_n68), .A(REG61_n83), .ZN(
        REG61_n55) );
  NAND2_X1 REG61_U20 ( .A1(temp6[5]), .A2(REG61_n43), .ZN(REG61_n84) );
  OAI21_X1 REG61_U19 ( .B1(REG61_n44), .B2(REG61_n67), .A(REG61_n84), .ZN(
        REG61_n56) );
  NAND2_X1 REG61_U18 ( .A1(temp6[1]), .A2(REG61_n43), .ZN(REG61_n88) );
  OAI21_X1 REG61_U17 ( .B1(REG61_n44), .B2(REG61_n63), .A(REG61_n88), .ZN(
        REG61_n60) );
  NAND2_X1 REG61_U16 ( .A1(temp6[0]), .A2(REG61_n43), .ZN(REG61_n89) );
  OAI21_X1 REG61_U15 ( .B1(REG61_n44), .B2(REG61_n62), .A(REG61_n89), .ZN(
        REG61_n61) );
  NAND2_X1 REG61_U14 ( .A1(temp6[11]), .A2(REG61_n43), .ZN(REG61_n78) );
  OAI21_X1 REG61_U13 ( .B1(REG61_n44), .B2(REG61_n73), .A(REG61_n78), .ZN(
        REG61_n50) );
  NAND2_X1 REG61_U12 ( .A1(temp6[12]), .A2(REG61_n43), .ZN(REG61_n77) );
  OAI21_X1 REG61_U11 ( .B1(REG61_n44), .B2(REG61_n74), .A(REG61_n77), .ZN(
        REG61_n49) );
  NAND2_X1 REG61_U10 ( .A1(temp6[10]), .A2(REG61_n44), .ZN(REG61_n79) );
  OAI21_X1 REG61_U9 ( .B1(REG61_n44), .B2(REG61_n72), .A(REG61_n79), .ZN(
        REG61_n51) );
  NAND2_X1 REG61_U8 ( .A1(temp6[13]), .A2(REG61_n43), .ZN(REG61_n76) );
  OAI21_X1 REG61_U7 ( .B1(REG61_n44), .B2(REG61_n75), .A(REG61_n76), .ZN(
        REG61_n48) );
  BUF_X1 REG61_U6 ( .A(n48), .Z(REG61_n47) );
  BUF_X1 REG61_U5 ( .A(n48), .Z(REG61_n46) );
  BUF_X1 REG61_U4 ( .A(VIN), .Z(REG61_n45) );
  BUF_X1 REG61_U3 ( .A(VIN), .Z(REG61_n43) );
  BUF_X1 REG61_U2 ( .A(VIN), .Z(REG61_n44) );
  DFFR_X1 REG61_q_reg_0_ ( .D(REG61_n61), .CK(CLK), .RN(REG61_n47), .Q(reg7[0]), .QN(REG61_n62) );
  DFFR_X1 REG61_q_reg_1_ ( .D(REG61_n60), .CK(CLK), .RN(REG61_n47), .Q(reg7[1]), .QN(REG61_n63) );
  DFFR_X1 REG61_q_reg_2_ ( .D(REG61_n59), .CK(CLK), .RN(REG61_n46), .Q(reg7[2]), .QN(REG61_n64) );
  DFFR_X1 REG61_q_reg_3_ ( .D(REG61_n58), .CK(CLK), .RN(REG61_n46), .Q(reg7[3]), .QN(REG61_n65) );
  DFFR_X1 REG61_q_reg_4_ ( .D(REG61_n57), .CK(CLK), .RN(REG61_n46), .Q(reg7[4]), .QN(REG61_n66) );
  DFFR_X1 REG61_q_reg_5_ ( .D(REG61_n56), .CK(CLK), .RN(REG61_n46), .Q(reg7[5]), .QN(REG61_n67) );
  DFFR_X1 REG61_q_reg_6_ ( .D(REG61_n55), .CK(CLK), .RN(REG61_n46), .Q(reg7[6]), .QN(REG61_n68) );
  DFFR_X1 REG61_q_reg_7_ ( .D(REG61_n54), .CK(CLK), .RN(REG61_n46), .Q(reg7[7]), .QN(REG61_n69) );
  DFFR_X1 REG61_q_reg_8_ ( .D(REG61_n53), .CK(CLK), .RN(REG61_n46), .Q(reg7[8]), .QN(REG61_n70) );
  DFFR_X1 REG61_q_reg_9_ ( .D(REG61_n52), .CK(CLK), .RN(REG61_n46), .Q(reg7[9]), .QN(REG61_n71) );
  DFFR_X1 REG61_q_reg_10_ ( .D(REG61_n51), .CK(CLK), .RN(REG61_n46), .Q(
        reg7[10]), .QN(REG61_n72) );
  DFFR_X1 REG61_q_reg_11_ ( .D(REG61_n50), .CK(CLK), .RN(REG61_n46), .Q(
        reg7[11]), .QN(REG61_n73) );
  DFFR_X1 REG61_q_reg_12_ ( .D(REG61_n49), .CK(CLK), .RN(REG61_n46), .Q(
        reg7[12]), .QN(REG61_n74) );
  DFFR_X1 REG61_q_reg_13_ ( .D(REG61_n48), .CK(CLK), .RN(REG61_n46), .Q(
        reg7[13]), .QN(REG61_n75) );
endmodule

