
module IIR_ADV ( CLK, RST_n, VIN, DIN, B0, B1, B2, B3, A1, A2, VOUT, DOUT );
  input [13:0] DIN;
  input [13:0] B0;
  input [13:0] B1;
  input [13:0] B2;
  input [13:0] B3;
  input [13:0] A1;
  input [13:0] A2;
  output [13:0] DOUT;
  input CLK, RST_n, VIN;
  output VOUT;
  wire   p6_final_product2_25_, p6_final_product2_26_, p6_muxs_out_3__6_,
         p6_muxs_out_3__7_, p6_muxs_out_3__8_, p6_muxs_out_3__9_,
         p6_muxs_out_3__10_, p6_muxs_out_3__11_, p6_muxs_out_3__12_,
         p6_muxs_out_3__13_, p6_muxs_out_3__14_, p6_muxs_out_3__15_,
         p6_muxs_out_3__16_, p6_muxs_out_3__17_, p6_muxs_out_3__18_,
         p6_muxs_out_3__19_, p6_muxs_out_3__20_, p6_muxs_out_2__6_,
         p6_muxs_out_2__7_, p6_muxs_out_2__8_, p6_muxs_out_2__9_,
         p6_muxs_out_2__10_, p6_muxs_out_2__11_, p6_muxs_out_2__12_,
         p6_muxs_out_2__13_, p6_muxs_out_2__14_, p6_muxs_out_2__15_,
         p6_muxs_out_2__16_, p6_muxs_out_2__17_, p6_muxs_out_2__18_,
         p6_muxs_out_1__6_, p6_muxs_out_1__8_, p6_muxs_out_1__9_,
         p6_muxs_out_1__10_, p6_muxs_out_1__11_, p6_muxs_out_1__12_,
         p6_muxs_out_1__13_, p6_muxs_out_1__14_, p6_muxs_out_1__15_,
         p6_muxs_out_1__16_, p6_minus_A_shifted_13_, p6_minus_A_shifted_14_,
         p6_minus_A_shifted_15_, p6_minus_A_shifted_16_,
         p6_minus_A_shifted_17_, p6_minus_A_shifted_18_,
         p6_minus_A_shifted_19_, p6_minus_A_shifted_20_,
         p6_minus_A_shifted_21_, p6_minus_A_shifted_22_,
         p6_minus_A_shifted_23_, p6_minus_A_shifted_25_,
         p6_minus_A_shifted_38_, p7_final_product2_25_, p7_final_product2_26_,
         p7_muxs_out_3__6_, p7_muxs_out_3__7_, p7_muxs_out_3__8_,
         p7_muxs_out_3__9_, p7_muxs_out_3__10_, p7_muxs_out_3__11_,
         p7_muxs_out_3__12_, p7_muxs_out_3__13_, p7_muxs_out_3__14_,
         p7_muxs_out_3__15_, p7_muxs_out_3__16_, p7_muxs_out_3__17_,
         p7_muxs_out_3__18_, p7_muxs_out_3__19_, p7_muxs_out_3__20_,
         p7_muxs_out_2__6_, p7_muxs_out_2__7_, p7_muxs_out_2__8_,
         p7_muxs_out_2__9_, p7_muxs_out_2__10_, p7_muxs_out_2__11_,
         p7_muxs_out_2__12_, p7_muxs_out_2__13_, p7_muxs_out_2__14_,
         p7_muxs_out_2__15_, p7_muxs_out_2__16_, p7_muxs_out_2__17_,
         p7_muxs_out_2__18_, p7_muxs_out_1__6_, p7_muxs_out_1__8_,
         p7_muxs_out_1__9_, p7_muxs_out_1__10_, p7_muxs_out_1__11_,
         p7_muxs_out_1__12_, p7_muxs_out_1__13_, p7_muxs_out_1__14_,
         p7_muxs_out_1__15_, p7_muxs_out_1__16_, p7_minus_A_shifted_13_,
         p7_minus_A_shifted_14_, p7_minus_A_shifted_15_,
         p7_minus_A_shifted_16_, p7_minus_A_shifted_17_,
         p7_minus_A_shifted_18_, p7_minus_A_shifted_19_,
         p7_minus_A_shifted_20_, p7_minus_A_shifted_21_,
         p7_minus_A_shifted_22_, p7_minus_A_shifted_23_,
         p7_minus_A_shifted_25_, p7_minus_A_shifted_38_, p8_final_product2_25_,
         p8_final_product2_26_, p8_muxs_out_3__6_, p8_muxs_out_3__7_,
         p8_muxs_out_3__8_, p8_muxs_out_3__9_, p8_muxs_out_3__10_,
         p8_muxs_out_3__11_, p8_muxs_out_3__12_, p8_muxs_out_3__13_,
         p8_muxs_out_3__14_, p8_muxs_out_3__15_, p8_muxs_out_3__16_,
         p8_muxs_out_3__17_, p8_muxs_out_3__18_, p8_muxs_out_3__19_,
         p8_muxs_out_3__20_, p8_muxs_out_2__6_, p8_muxs_out_2__7_,
         p8_muxs_out_2__8_, p8_muxs_out_2__9_, p8_muxs_out_2__10_,
         p8_muxs_out_2__11_, p8_muxs_out_2__12_, p8_muxs_out_2__13_,
         p8_muxs_out_2__14_, p8_muxs_out_2__15_, p8_muxs_out_2__16_,
         p8_muxs_out_2__17_, p8_muxs_out_2__18_, p8_muxs_out_1__6_,
         p8_muxs_out_1__8_, p8_muxs_out_1__9_, p8_muxs_out_1__10_,
         p8_muxs_out_1__11_, p8_muxs_out_1__12_, p8_muxs_out_1__13_,
         p8_muxs_out_1__14_, p8_muxs_out_1__15_, p8_muxs_out_1__16_,
         p8_minus_A_shifted_13_, p8_minus_A_shifted_14_,
         p8_minus_A_shifted_15_, p8_minus_A_shifted_16_,
         p8_minus_A_shifted_17_, p8_minus_A_shifted_18_,
         p8_minus_A_shifted_19_, p8_minus_A_shifted_20_,
         p8_minus_A_shifted_21_, p8_minus_A_shifted_22_,
         p8_minus_A_shifted_23_, p8_minus_A_shifted_25_,
         p8_minus_A_shifted_38_, p9_final_product2_25_, p9_final_product2_26_,
         p9_muxs_out_3__6_, p9_muxs_out_3__7_, p9_muxs_out_3__8_,
         p9_muxs_out_3__9_, p9_muxs_out_3__10_, p9_muxs_out_3__11_,
         p9_muxs_out_3__12_, p9_muxs_out_3__13_, p9_muxs_out_3__14_,
         p9_muxs_out_3__15_, p9_muxs_out_3__16_, p9_muxs_out_3__17_,
         p9_muxs_out_3__18_, p9_muxs_out_3__19_, p9_muxs_out_3__20_,
         p9_muxs_out_2__6_, p9_muxs_out_2__7_, p9_muxs_out_2__8_,
         p9_muxs_out_2__9_, p9_muxs_out_2__10_, p9_muxs_out_2__11_,
         p9_muxs_out_2__12_, p9_muxs_out_2__13_, p9_muxs_out_2__14_,
         p9_muxs_out_2__15_, p9_muxs_out_2__16_, p9_muxs_out_2__17_,
         p9_muxs_out_2__18_, p9_muxs_out_1__6_, p9_muxs_out_1__8_,
         p9_muxs_out_1__9_, p9_muxs_out_1__10_, p9_muxs_out_1__11_,
         p9_muxs_out_1__12_, p9_muxs_out_1__13_, p9_muxs_out_1__14_,
         p9_muxs_out_1__15_, p9_muxs_out_1__16_, p9_minus_A_shifted_13_,
         p9_minus_A_shifted_14_, p9_minus_A_shifted_15_,
         p9_minus_A_shifted_16_, p9_minus_A_shifted_17_,
         p9_minus_A_shifted_18_, p9_minus_A_shifted_19_,
         p9_minus_A_shifted_20_, p9_minus_A_shifted_21_,
         p9_minus_A_shifted_22_, p9_minus_A_shifted_23_,
         p9_minus_A_shifted_25_, p9_minus_A_shifted_38_,
         p11_final_product2_25_, p11_final_product2_26_, p11_muxs_out_3__6_,
         p11_muxs_out_3__7_, p11_muxs_out_3__8_, p11_muxs_out_3__9_,
         p11_muxs_out_3__10_, p11_muxs_out_3__11_, p11_muxs_out_3__12_,
         p11_muxs_out_3__13_, p11_muxs_out_3__14_, p11_muxs_out_3__15_,
         p11_muxs_out_3__16_, p11_muxs_out_3__17_, p11_muxs_out_3__18_,
         p11_muxs_out_3__19_, p11_muxs_out_3__20_, p11_muxs_out_2__6_,
         p11_muxs_out_2__7_, p11_muxs_out_2__8_, p11_muxs_out_2__9_,
         p11_muxs_out_2__10_, p11_muxs_out_2__11_, p11_muxs_out_2__12_,
         p11_muxs_out_2__13_, p11_muxs_out_2__14_, p11_muxs_out_2__15_,
         p11_muxs_out_2__16_, p11_muxs_out_2__17_, p11_muxs_out_2__18_,
         p11_muxs_out_1__6_, p11_muxs_out_1__8_, p11_muxs_out_1__9_,
         p11_muxs_out_1__10_, p11_muxs_out_1__11_, p11_muxs_out_1__12_,
         p11_muxs_out_1__13_, p11_muxs_out_1__14_, p11_muxs_out_1__15_,
         p11_muxs_out_1__16_, p11_minus_A_shifted_14_, p11_minus_A_shifted_16_,
         p10_final_product2_25_, p10_final_product2_26_, p10_muxs_out_3__6_,
         p10_muxs_out_3__7_, p10_muxs_out_3__8_, p10_muxs_out_3__9_,
         p10_muxs_out_3__10_, p10_muxs_out_3__11_, p10_muxs_out_3__12_,
         p10_muxs_out_3__13_, p10_muxs_out_3__14_, p10_muxs_out_3__15_,
         p10_muxs_out_3__16_, p10_muxs_out_3__17_, p10_muxs_out_3__18_,
         p10_muxs_out_3__19_, p10_muxs_out_3__20_, p10_muxs_out_2__6_,
         p10_muxs_out_2__7_, p10_muxs_out_2__8_, p10_muxs_out_2__9_,
         p10_muxs_out_2__10_, p10_muxs_out_2__11_, p10_muxs_out_2__12_,
         p10_muxs_out_2__13_, p10_muxs_out_2__14_, p10_muxs_out_2__15_,
         p10_muxs_out_2__16_, p10_muxs_out_2__17_, p10_muxs_out_2__18_,
         p10_muxs_out_1__6_, p10_muxs_out_1__8_, p10_muxs_out_1__9_,
         p10_muxs_out_1__10_, p10_muxs_out_1__11_, p10_muxs_out_1__12_,
         p10_muxs_out_1__13_, p10_muxs_out_1__14_, p10_muxs_out_1__15_,
         p10_muxs_out_1__16_, p10_minus_A_shifted_14_, p10_minus_A_shifted_16_,
         n14, n15, n16, n17, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n275, n276, n277, n278, n279,
         n280, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n336,
         n337, n338, n339, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n601, n602, n603, n604, n605, n606,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n662, n663,
         n664, n665, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n927, n928, n929, n930, n931, n932, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n988, n989, n990,
         n991, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1253, n1254, n1255, n1256,
         n1257, n1258, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1314, n1315, n1316, n1317, n1319,
         n1321, n1322, n1323, n1324, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1402, n1403,
         n1404, n1405, n1406, n1407, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1447,
         n1448, n1449, n1450, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1554, n1555, n1556, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1653, n1654, n1655, n1656, n1657, n1658,
         n1660, n1661, n1662, n1663, n1665, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1742, n1743,
         n1744, n1745, n1746, n1747, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1787,
         n1788, n1789, n1790, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1894, n1895, n1896, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2074,
         n2077, n2083, n2087, n2093, n2100, n2104, n2107, n2110, n2113, n2116,
         n2117, n2118, n2119, n2120, n2122, n2125, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, s8_add_23_DP_OP_277_3998_2_n91,
         s8_add_23_DP_OP_277_3998_2_n90, s8_add_23_DP_OP_277_3998_2_n89,
         s8_add_23_DP_OP_277_3998_2_n88, s8_add_23_DP_OP_277_3998_2_n87,
         s8_add_23_DP_OP_277_3998_2_n86, s8_add_23_DP_OP_277_3998_2_n85,
         s8_add_23_DP_OP_277_3998_2_n84, s8_add_23_DP_OP_277_3998_2_n83,
         s8_add_23_DP_OP_277_3998_2_n82, s8_add_23_DP_OP_277_3998_2_n81,
         s8_add_23_DP_OP_277_3998_2_n80, s8_add_23_DP_OP_277_3998_2_n79,
         s8_add_23_DP_OP_277_3998_2_n78, s8_add_23_DP_OP_277_3998_2_n77,
         s8_add_23_DP_OP_277_3998_2_n76, s8_add_23_DP_OP_277_3998_2_n75,
         s8_add_23_DP_OP_277_3998_2_n74, s8_add_23_DP_OP_277_3998_2_n73,
         s8_add_23_DP_OP_277_3998_2_n72, s8_add_23_DP_OP_277_3998_2_n71,
         s8_add_23_DP_OP_277_3998_2_n70, s8_add_23_DP_OP_277_3998_2_n69,
         s8_add_23_DP_OP_277_3998_2_n68, s8_add_23_DP_OP_277_3998_2_n67,
         s8_add_23_DP_OP_277_3998_2_n66, s8_add_23_DP_OP_277_3998_2_n65,
         s8_add_23_DP_OP_277_3998_2_n64, s8_add_23_DP_OP_277_3998_2_n63,
         s8_add_23_DP_OP_277_3998_2_n62, s8_add_23_DP_OP_277_3998_2_n61,
         s8_add_23_DP_OP_277_3998_2_n60, s8_add_23_DP_OP_277_3998_2_n59,
         s8_add_23_DP_OP_277_3998_2_n58, s8_add_23_DP_OP_277_3998_2_n57,
         s8_add_23_DP_OP_277_3998_2_n56, s8_add_23_DP_OP_277_3998_2_n55,
         s8_add_23_DP_OP_277_3998_2_n54, s8_add_23_DP_OP_277_3998_2_n53,
         s8_add_23_DP_OP_277_3998_2_n52, s8_add_23_DP_OP_277_3998_2_n51,
         s8_add_23_DP_OP_277_3998_2_n50, s8_add_23_DP_OP_277_3998_2_n49,
         s8_add_23_DP_OP_277_3998_2_n48, s8_add_23_DP_OP_277_3998_2_n47,
         s8_add_23_DP_OP_277_3998_2_n46, s8_add_23_DP_OP_277_3998_2_n45,
         s8_add_23_DP_OP_277_3998_2_n44, s8_add_23_DP_OP_277_3998_2_n43,
         s8_add_23_DP_OP_277_3998_2_n42, s8_add_23_DP_OP_277_3998_2_n39,
         s8_add_23_DP_OP_277_3998_2_n38, s8_add_23_DP_OP_277_3998_2_n37,
         s8_add_23_DP_OP_277_3998_2_n36, s8_add_23_DP_OP_277_3998_2_n35,
         s8_add_23_DP_OP_277_3998_2_n34, s8_add_23_DP_OP_277_3998_2_n33,
         s8_add_23_DP_OP_277_3998_2_n32, s8_add_23_DP_OP_277_3998_2_n31,
         s8_add_23_DP_OP_277_3998_2_n30, s8_add_23_DP_OP_277_3998_2_n29,
         s8_add_23_DP_OP_277_3998_2_n28, s8_add_23_DP_OP_277_3998_2_n27,
         s9_add_23_DP_OP_276_9387_1_n60, s9_add_23_DP_OP_276_9387_1_n59,
         s9_add_23_DP_OP_276_9387_1_n58, s9_add_23_DP_OP_276_9387_1_n57,
         s9_add_23_DP_OP_276_9387_1_n56, s9_add_23_DP_OP_276_9387_1_n55,
         s9_add_23_DP_OP_276_9387_1_n54, s9_add_23_DP_OP_276_9387_1_n53,
         s9_add_23_DP_OP_276_9387_1_n52, s9_add_23_DP_OP_276_9387_1_n51,
         s9_add_23_DP_OP_276_9387_1_n50, s9_add_23_DP_OP_276_9387_1_n49,
         s9_add_23_DP_OP_276_9387_1_n48, s9_add_23_DP_OP_276_9387_1_n47,
         s9_add_23_DP_OP_276_9387_1_n46, s9_add_23_DP_OP_276_9387_1_n45,
         s9_add_23_DP_OP_276_9387_1_n44, s9_add_23_DP_OP_276_9387_1_n43,
         s9_add_23_DP_OP_276_9387_1_n42, s9_add_23_DP_OP_276_9387_1_n41,
         s9_add_23_DP_OP_276_9387_1_n40, s9_add_23_DP_OP_276_9387_1_n39,
         s9_add_23_DP_OP_276_9387_1_n38, s9_add_23_DP_OP_276_9387_1_n37,
         s9_add_23_DP_OP_276_9387_1_n34, s9_add_23_DP_OP_276_9387_1_n33,
         s9_add_23_DP_OP_276_9387_1_n32, s9_add_23_DP_OP_276_9387_1_n31,
         s9_add_23_DP_OP_276_9387_1_n30, s9_add_23_DP_OP_276_9387_1_n29,
         s9_add_23_DP_OP_276_9387_1_n28, s9_add_23_DP_OP_276_9387_1_n27,
         s9_add_23_DP_OP_276_9387_1_n26, s9_add_23_DP_OP_276_9387_1_n25,
         s9_add_23_DP_OP_276_9387_1_n24, s9_add_23_DP_OP_276_9387_1_n23,
         s9_add_23_DP_OP_276_9387_1_n22,
         p10_Partial_products_sum_add_23_carry_7_,
         p10_Partial_products_sum_add_23_carry_8_,
         p10_Partial_products_sum_add_23_carry_9_,
         p10_Partial_products_sum_add_23_carry_10_,
         p10_Partial_products_sum_add_23_carry_11_,
         p10_Partial_products_sum_add_23_carry_12_,
         p10_Partial_products_sum_add_23_carry_13_,
         p10_Partial_products_sum_add_23_carry_14_,
         p10_Partial_products_sum_add_23_carry_15_,
         p10_Partial_products_sum_add_23_carry_16_,
         p10_Partial_products_sum_add_23_carry_17_,
         p10_Partial_products_sum_add_23_carry_18_,
         p10_Partial_products_sum_add_23_carry_19_,
         p10_Partial_products_sum_add_23_carry_20_,
         p11_Partial_products_sum_add_23_carry_7_,
         p11_Partial_products_sum_add_23_carry_8_,
         p11_Partial_products_sum_add_23_carry_9_,
         p11_Partial_products_sum_add_23_carry_10_,
         p11_Partial_products_sum_add_23_carry_11_,
         p11_Partial_products_sum_add_23_carry_12_,
         p11_Partial_products_sum_add_23_carry_13_,
         p11_Partial_products_sum_add_23_carry_14_,
         p11_Partial_products_sum_add_23_carry_15_,
         p11_Partial_products_sum_add_23_carry_16_,
         p11_Partial_products_sum_add_23_carry_17_,
         p11_Partial_products_sum_add_23_carry_18_,
         p11_Partial_products_sum_add_23_carry_19_,
         p11_Partial_products_sum_add_23_carry_20_,
         p9_Partial_products_sum_add_23_carry_7_,
         p9_Partial_products_sum_add_23_carry_8_,
         p9_Partial_products_sum_add_23_carry_9_,
         p9_Partial_products_sum_add_23_carry_10_,
         p9_Partial_products_sum_add_23_carry_11_,
         p9_Partial_products_sum_add_23_carry_12_,
         p9_Partial_products_sum_add_23_carry_13_,
         p9_Partial_products_sum_add_23_carry_14_,
         p9_Partial_products_sum_add_23_carry_15_,
         p9_Partial_products_sum_add_23_carry_16_,
         p9_Partial_products_sum_add_23_carry_17_,
         p9_Partial_products_sum_add_23_carry_18_,
         p9_Partial_products_sum_add_23_carry_19_,
         p9_Partial_products_sum_add_23_carry_20_,
         p9_Partial_products_sum_add_23_B_0_,
         p8_Partial_products_sum_add_23_carry_7_,
         p8_Partial_products_sum_add_23_carry_8_,
         p8_Partial_products_sum_add_23_carry_9_,
         p8_Partial_products_sum_add_23_carry_10_,
         p8_Partial_products_sum_add_23_carry_11_,
         p8_Partial_products_sum_add_23_carry_12_,
         p8_Partial_products_sum_add_23_carry_13_,
         p8_Partial_products_sum_add_23_carry_14_,
         p8_Partial_products_sum_add_23_carry_15_,
         p8_Partial_products_sum_add_23_carry_16_,
         p8_Partial_products_sum_add_23_carry_17_,
         p8_Partial_products_sum_add_23_carry_18_,
         p8_Partial_products_sum_add_23_carry_19_,
         p8_Partial_products_sum_add_23_carry_20_,
         p8_Partial_products_sum_add_23_B_0_,
         p7_Partial_products_sum_add_23_carry_7_,
         p7_Partial_products_sum_add_23_carry_8_,
         p7_Partial_products_sum_add_23_carry_9_,
         p7_Partial_products_sum_add_23_carry_10_,
         p7_Partial_products_sum_add_23_carry_11_,
         p7_Partial_products_sum_add_23_carry_12_,
         p7_Partial_products_sum_add_23_carry_13_,
         p7_Partial_products_sum_add_23_carry_14_,
         p7_Partial_products_sum_add_23_carry_15_,
         p7_Partial_products_sum_add_23_carry_16_,
         p7_Partial_products_sum_add_23_carry_17_,
         p7_Partial_products_sum_add_23_carry_18_,
         p7_Partial_products_sum_add_23_carry_19_,
         p7_Partial_products_sum_add_23_carry_20_,
         p7_Partial_products_sum_add_23_B_0_,
         p6_Partial_products_sum_add_23_B_0_,
         p6_Partial_products_sum_add_23_n15,
         p6_Partial_products_sum_add_23_n14,
         p6_Partial_products_sum_add_23_n13,
         p6_Partial_products_sum_add_23_n12,
         p6_Partial_products_sum_add_23_n11,
         p6_Partial_products_sum_add_23_n10, p6_Partial_products_sum_add_23_n9,
         p6_Partial_products_sum_add_23_n8, p6_Partial_products_sum_add_23_n7,
         p6_Partial_products_sum_add_23_n6, p6_Partial_products_sum_add_23_n5,
         p6_Partial_products_sum_add_23_n4, p6_Partial_products_sum_add_23_n3,
         p6_Partial_products_sum_add_23_n2, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440;
  wire   [13:0] xin;
  wire   [13:0] w;
  wire   [13:0] reg1_reg;
  wire   [13:0] temp1;
  wire   [13:0] mul1_reg;
  wire   [13:0] reg2;
  wire   [13:0] reg2_reg;
  wire   [13:0] temp2;
  wire   [13:0] mul2_reg;
  wire   [13:0] reg3_reg;
  wire   [13:0] temp3;
  wire   [13:0] mul3_reg;
  wire   [13:0] reg4_reg;
  wire   [13:0] temp4;
  wire   [13:0] mul4_reg;
  wire   [13:0] temp6;
  wire   [13:0] reg4;
  wire   [13:0] temp5;
  wire   [13:0] reg6;
  wire   [13:0] reg7;
  wire   [13:0] ff;
  wire   [72:54] p6_C;
  wire   [72:54] p6_S;
  wire   [26:26] p7_final_product1;
  wire   [72:54] p7_C;
  wire   [72:54] p7_S;
  wire   [26:26] p8_final_product1;
  wire   [72:54] p8_C;
  wire   [72:54] p8_S;
  wire   [26:26] p9_final_product1;
  wire   [72:54] p9_C;
  wire   [72:54] p9_S;
  wire   [26:26] p11_final_product1;
  wire   [72:54] p11_C;
  wire   [72:54] p11_S;
  wire   [26:26] p10_final_product1;
  wire   [72:54] p10_C;
  wire   [72:54] p10_S;

  DFFR_X1 xin_in_reg_13_ ( .D(n2595), .CK(CLK), .RN(RST_n), .Q(n2240) );
  DFFR_X1 xin_in_reg_12_ ( .D(n2594), .CK(CLK), .RN(RST_n), .Q(n2239) );
  DFFR_X1 xin_in_reg_11_ ( .D(n2593), .CK(CLK), .RN(RST_n), .Q(n2238) );
  DFFR_X1 xin_in_reg_10_ ( .D(n2592), .CK(CLK), .RN(RST_n), .Q(n2237) );
  DFFR_X1 xin_in_reg_9_ ( .D(n2591), .CK(CLK), .RN(RST_n), .Q(n2236) );
  DFFR_X1 xin_in_reg_8_ ( .D(n2590), .CK(CLK), .RN(RST_n), .Q(n2235) );
  DFFR_X1 xin_in_reg_7_ ( .D(n2589), .CK(CLK), .RN(RST_n), .Q(n2234) );
  DFFR_X1 xin_in_reg_6_ ( .D(n2588), .CK(CLK), .RN(RST_n), .Q(n2233) );
  DFFR_X1 xin_in_reg_5_ ( .D(n2587), .CK(CLK), .RN(RST_n), .Q(n2232) );
  DFFR_X1 xin_in_reg_4_ ( .D(n2586), .CK(CLK), .RN(RST_n), .Q(n2231) );
  DFFR_X1 xin_in_reg_3_ ( .D(n2585), .CK(CLK), .RN(RST_n), .Q(n2230) );
  DFFR_X1 xin_in_reg_2_ ( .D(n2584), .CK(CLK), .RN(RST_n), .Q(n2229) );
  DFFR_X1 xin_in_reg_1_ ( .D(n2583), .CK(CLK), .RN(RST_n), .Q(n2228) );
  DFFR_X1 xin_in_reg_0_ ( .D(n2582), .CK(CLK), .RN(RST_n), .Q(n2227) );
  DFFR_X1 VOUT_reg ( .D(n2581), .CK(CLK), .RN(RST_n), .Q(VOUT), .QN(n2226) );
  DFFR_X1 REGISTER_in_q_reg_0_ ( .D(n2580), .CK(CLK), .RN(RST_n), .Q(xin[0])
         );
  DFFR_X1 REGISTER_in_q_reg_1_ ( .D(n2579), .CK(CLK), .RN(RST_n), .Q(xin[1]), 
        .QN(n2682) );
  DFFR_X1 REGISTER_in_q_reg_2_ ( .D(n2578), .CK(CLK), .RN(RST_n), .Q(xin[2])
         );
  DFFR_X1 REGISTER_in_q_reg_3_ ( .D(n2577), .CK(CLK), .RN(RST_n), .Q(xin[3])
         );
  DFFR_X1 REGISTER_in_q_reg_4_ ( .D(n2576), .CK(CLK), .RN(RST_n), .Q(xin[4])
         );
  DFFR_X1 REGISTER_in_q_reg_5_ ( .D(n2575), .CK(CLK), .RN(RST_n), .Q(xin[5])
         );
  DFFR_X1 REGISTER_in_q_reg_6_ ( .D(n2574), .CK(CLK), .RN(RST_n), .Q(xin[6])
         );
  DFFR_X1 REGISTER_in_q_reg_7_ ( .D(n2573), .CK(CLK), .RN(RST_n), .Q(xin[7])
         );
  DFFR_X1 REGISTER_in_q_reg_8_ ( .D(n2572), .CK(CLK), .RN(RST_n), .Q(xin[8])
         );
  DFFR_X1 REGISTER_in_q_reg_9_ ( .D(n2571), .CK(CLK), .RN(RST_n), .Q(xin[9])
         );
  DFFR_X1 REGISTER_in_q_reg_10_ ( .D(n2570), .CK(CLK), .RN(RST_n), .Q(xin[10])
         );
  DFFR_X1 REGISTER_in_q_reg_11_ ( .D(n2569), .CK(CLK), .RN(RST_n), .Q(xin[11])
         );
  DFFR_X1 REGISTER_in_q_reg_12_ ( .D(n2568), .CK(CLK), .RN(RST_n), .Q(xin[12])
         );
  DFFR_X1 REGISTER_in_q_reg_13_ ( .D(n2567), .CK(CLK), .RN(RST_n), .Q(xin[13])
         );
  DFFR_X1 REG61_q_reg_13_ ( .D(n2566), .CK(CLK), .RN(RST_n), .Q(reg7[13]) );
  DFFR_X1 REGISTER1_q_reg_0_ ( .D(n2565), .CK(CLK), .RN(RST_n), .Q(reg1_reg[0]), .QN(n2836) );
  DFFR_X1 REG11_q_reg_0_ ( .D(n2564), .CK(CLK), .RN(RST_n), .Q(reg2[0]), .QN(
        n2838) );
  DFFR_X1 REGISTER2_q_reg_0_ ( .D(n2563), .CK(CLK), .RN(RST_n), .Q(reg2_reg[0]), .QN(n2837) );
  DFFR_X1 REG21_q_reg_0_ ( .D(n2562), .CK(CLK), .RN(RST_n), .QN(n2868) );
  DFFR_X1 REGISTER3_q_reg_0_ ( .D(n2561), .CK(CLK), .RN(RST_n), .Q(reg3_reg[0]), .QN(n2797) );
  DFFR_X1 REG31_q_reg_0_ ( .D(n2560), .CK(CLK), .RN(RST_n), .Q(reg4[0]), .QN(
        n2839) );
  DFFR_X1 REG41_q_reg_0_ ( .D(n2559), .CK(CLK), .RN(RST_n), .QN(n2869) );
  DFFR_X1 REGISTER4_q_reg_0_ ( .D(n2558), .CK(CLK), .RN(RST_n), .Q(reg4_reg[0]), .QN(n2798) );
  DFFR_X1 REGISTER1_q_reg_1_ ( .D(n2557), .CK(CLK), .RN(RST_n), .Q(reg1_reg[1]), .QN(n2864) );
  DFFR_X1 REG11_q_reg_1_ ( .D(n2556), .CK(CLK), .RN(RST_n), .Q(reg2[1]), .QN(
        p11_minus_A_shifted_14_) );
  DFFR_X1 REGISTER2_q_reg_1_ ( .D(n2555), .CK(CLK), .RN(RST_n), .Q(reg2_reg[1]), .QN(n2865) );
  DFFR_X1 REG21_q_reg_1_ ( .D(n2554), .CK(CLK), .RN(RST_n), .Q(n2223) );
  DFFR_X1 REGISTER3_q_reg_1_ ( .D(n2553), .CK(CLK), .RN(RST_n), .Q(reg3_reg[1]), .QN(n2840) );
  DFFR_X1 REG31_q_reg_1_ ( .D(n2552), .CK(CLK), .RN(RST_n), .Q(reg4[1]), .QN(
        p10_minus_A_shifted_14_) );
  DFFR_X1 REG41_q_reg_1_ ( .D(n2551), .CK(CLK), .RN(RST_n), .Q(n2222) );
  DFFR_X1 REGISTER4_q_reg_1_ ( .D(n2550), .CK(CLK), .RN(RST_n), .Q(reg4_reg[1]), .QN(n2841) );
  DFFR_X1 REGISTER1_q_reg_2_ ( .D(n2549), .CK(CLK), .RN(RST_n), .Q(reg1_reg[2]), .QN(n2792) );
  DFFR_X1 REG11_q_reg_2_ ( .D(n2548), .CK(CLK), .RN(RST_n), .Q(reg2[2]), .QN(
        n2820) );
  DFFR_X1 REGISTER2_q_reg_2_ ( .D(n2547), .CK(CLK), .RN(RST_n), .Q(reg2_reg[2]), .QN(n2793) );
  DFFR_X1 REG21_q_reg_2_ ( .D(n2546), .CK(CLK), .RN(RST_n), .Q(n2221), .QN(
        n2888) );
  DFFR_X1 REGISTER3_q_reg_2_ ( .D(n2545), .CK(CLK), .RN(RST_n), .Q(reg3_reg[2]), .QN(n2794) );
  DFFR_X1 REG31_q_reg_2_ ( .D(n2544), .CK(CLK), .RN(RST_n), .Q(reg4[2]), .QN(
        n2821) );
  DFFR_X1 REG41_q_reg_2_ ( .D(n2543), .CK(CLK), .RN(RST_n), .Q(n2220), .QN(
        n2889) );
  DFFR_X1 REGISTER4_q_reg_2_ ( .D(n2542), .CK(CLK), .RN(RST_n), .Q(reg4_reg[2]), .QN(n2795) );
  DFFR_X1 REG11_q_reg_3_ ( .D(n2540), .CK(CLK), .RN(RST_n), .Q(reg2[3]), .QN(
        p11_minus_A_shifted_16_) );
  DFFR_X1 REG21_q_reg_3_ ( .D(n2538), .CK(CLK), .RN(RST_n), .Q(n2219), .QN(
        n2890) );
  DFFR_X1 REG31_q_reg_3_ ( .D(n2536), .CK(CLK), .RN(RST_n), .Q(reg4[3]), .QN(
        p10_minus_A_shifted_16_) );
  DFFR_X1 REG41_q_reg_3_ ( .D(n2535), .CK(CLK), .RN(RST_n), .Q(n2218), .QN(
        n2891) );
  DFFR_X1 REG11_q_reg_4_ ( .D(n2532), .CK(CLK), .RN(RST_n), .Q(reg2[4]), .QN(
        n2817) );
  DFFR_X1 REGISTER2_q_reg_4_ ( .D(n2531), .CK(CLK), .RN(RST_n), .Q(reg2_reg[4]), .QN(n2827) );
  DFFR_X1 REG21_q_reg_4_ ( .D(n2530), .CK(CLK), .RN(RST_n), .Q(n2217), .QN(
        n2892) );
  DFFR_X1 REG31_q_reg_4_ ( .D(n2528), .CK(CLK), .RN(RST_n), .Q(reg4[4]), .QN(
        n2818) );
  DFFR_X1 REG41_q_reg_4_ ( .D(n2527), .CK(CLK), .RN(RST_n), .Q(n2216), .QN(
        n2893) );
  DFFR_X1 REG21_q_reg_5_ ( .D(n2522), .CK(CLK), .RN(RST_n), .Q(n2215), .QN(
        n2894) );
  DFFR_X1 REG31_q_reg_5_ ( .D(n2520), .CK(CLK), .RN(RST_n), .Q(reg4[5]), .QN(
        n2813) );
  DFFR_X1 REG41_q_reg_5_ ( .D(n2519), .CK(CLK), .RN(RST_n), .Q(n2214), .QN(
        n2895) );
  DFFR_X1 REG21_q_reg_6_ ( .D(n2514), .CK(CLK), .RN(RST_n), .Q(n2213), .QN(
        n2896) );
  DFFR_X1 REG31_q_reg_6_ ( .D(n2512), .CK(CLK), .RN(RST_n), .Q(reg4[6]), .QN(
        n2815) );
  DFFR_X1 REG41_q_reg_6_ ( .D(n2511), .CK(CLK), .RN(RST_n), .Q(n2212), .QN(
        n2897) );
  DFFR_X1 REG21_q_reg_7_ ( .D(n2506), .CK(CLK), .RN(RST_n), .QN(n2870) );
  DFFR_X1 REG41_q_reg_7_ ( .D(n2503), .CK(CLK), .RN(RST_n), .QN(n2871) );
  DFFR_X1 REGISTER1_q_reg_8_ ( .D(n2501), .CK(CLK), .RN(RST_n), .Q(reg1_reg[8]), .QN(n2881) );
  DFFR_X1 REG11_q_reg_8_ ( .D(n2500), .CK(CLK), .RN(RST_n), .Q(reg2[8]), .QN(
        n2811) );
  DFFR_X1 REGISTER2_q_reg_8_ ( .D(n2499), .CK(CLK), .RN(RST_n), .Q(reg2_reg[8]), .QN(n2885) );
  DFFR_X1 REG21_q_reg_8_ ( .D(n2498), .CK(CLK), .RN(RST_n), .QN(n2806) );
  DFFR_X1 REGISTER3_q_reg_8_ ( .D(n2497), .CK(CLK), .RN(RST_n), .Q(reg3_reg[8]), .QN(n2886) );
  DFFR_X1 REG41_q_reg_8_ ( .D(n2495), .CK(CLK), .RN(RST_n), .QN(n2807) );
  DFFR_X1 REGISTER4_q_reg_8_ ( .D(n2494), .CK(CLK), .RN(RST_n), .Q(reg4_reg[8]), .QN(n2887) );
  DFFR_X1 REGISTER1_q_reg_9_ ( .D(n2493), .CK(CLK), .RN(RST_n), .Q(reg1_reg[9]), .QN(n2819) );
  DFFR_X1 REG11_q_reg_9_ ( .D(n2492), .CK(CLK), .RN(RST_n), .Q(reg2[9]), .QN(
        n2816) );
  DFFR_X1 REGISTER2_q_reg_9_ ( .D(n2491), .CK(CLK), .RN(RST_n), .Q(reg2_reg[9]), .QN(n2812) );
  DFFR_X1 REG21_q_reg_9_ ( .D(n2490), .CK(CLK), .RN(RST_n), .QN(n2872) );
  DFFR_X1 REGISTER3_q_reg_9_ ( .D(n2489), .CK(CLK), .RN(RST_n), .Q(reg3_reg[9]), .QN(n2788) );
  DFFR_X1 REG31_q_reg_9_ ( .D(n2488), .CK(CLK), .RN(RST_n), .Q(reg4[9]), .QN(
        n2814) );
  DFFR_X1 REG41_q_reg_9_ ( .D(n2487), .CK(CLK), .RN(RST_n), .QN(n2873) );
  DFFR_X1 REGISTER4_q_reg_9_ ( .D(n2486), .CK(CLK), .RN(RST_n), .Q(reg4_reg[9]), .QN(n2789) );
  DFFR_X1 REGISTER1_q_reg_10_ ( .D(n2485), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[10]), .QN(n2880) );
  DFFR_X1 REGISTER2_q_reg_10_ ( .D(n2483), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[10]), .QN(n2882) );
  DFFR_X1 REG21_q_reg_10_ ( .D(n2482), .CK(CLK), .RN(RST_n), .QN(n2808) );
  DFFR_X1 REGISTER3_q_reg_10_ ( .D(n2481), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[10]), .QN(n2883) );
  DFFR_X1 REG31_q_reg_10_ ( .D(n2480), .CK(CLK), .RN(RST_n), .Q(reg4[10]), 
        .QN(n2810) );
  DFFR_X1 REG41_q_reg_10_ ( .D(n2479), .CK(CLK), .RN(RST_n), .QN(n2809) );
  DFFR_X1 REGISTER4_q_reg_10_ ( .D(n2478), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[10]), .QN(n2884) );
  DFFR_X1 REGISTER1_q_reg_11_ ( .D(n2477), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[11]), .QN(n2790) );
  DFFR_X1 REGISTER2_q_reg_11_ ( .D(n2475), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[11]), .QN(n2791) );
  DFFR_X1 REG21_q_reg_11_ ( .D(n2474), .CK(CLK), .RN(RST_n), .QN(n2874) );
  DFFR_X1 REGISTER3_q_reg_11_ ( .D(n2473), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[11]), .QN(n2786) );
  DFFR_X1 REG41_q_reg_11_ ( .D(n2471), .CK(CLK), .RN(RST_n), .QN(n2875) );
  DFFR_X1 REGISTER4_q_reg_11_ ( .D(n2470), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[11]), .QN(n2787) );
  DFFR_X1 REGISTER1_q_reg_12_ ( .D(n2469), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[12]), .QN(n2848) );
  DFFR_X1 REGISTER2_q_reg_12_ ( .D(n2467), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[12]), .QN(n2849) );
  DFFR_X1 REG21_q_reg_12_ ( .D(n2466), .CK(CLK), .RN(RST_n), .QN(n2876) );
  DFFR_X1 REGISTER3_q_reg_12_ ( .D(n2465), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[12]), .QN(n2802) );
  DFFR_X1 REG31_q_reg_12_ ( .D(n2464), .CK(CLK), .RN(RST_n), .Q(reg4[12]), 
        .QN(n2858) );
  DFFR_X1 REG41_q_reg_12_ ( .D(n2463), .CK(CLK), .RN(RST_n), .QN(n2877) );
  DFFR_X1 REGISTER4_q_reg_12_ ( .D(n2462), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[12]), .QN(n2803) );
  DFFR_X1 REGISTER1_q_reg_13_ ( .D(n2461), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[13]), .QN(n2867) );
  DFFR_X1 REG1_1_q_reg_0_ ( .D(n2460), .CK(CLK), .RN(RST_n), .Q(mul1_reg[0]), 
        .QN(n2199) );
  DFFR_X1 REG1_1_q_reg_1_ ( .D(n2459), .CK(CLK), .RN(RST_n), .Q(mul1_reg[1]), 
        .QN(n2198) );
  DFFR_X1 REG1_1_q_reg_2_ ( .D(n2458), .CK(CLK), .RN(RST_n), .Q(mul1_reg[2]), 
        .QN(n2197) );
  DFFR_X1 REG1_1_q_reg_3_ ( .D(n2457), .CK(CLK), .RN(RST_n), .Q(mul1_reg[3]), 
        .QN(n2196) );
  DFFR_X1 REG1_1_q_reg_4_ ( .D(n2456), .CK(CLK), .RN(RST_n), .Q(mul1_reg[4]), 
        .QN(n2195) );
  DFFR_X1 REG1_1_q_reg_5_ ( .D(n2455), .CK(CLK), .RN(RST_n), .Q(mul1_reg[5]), 
        .QN(n2194) );
  DFFR_X1 REG1_1_q_reg_6_ ( .D(n2454), .CK(CLK), .RN(RST_n), .Q(mul1_reg[6]), 
        .QN(n2193) );
  DFFR_X1 REG1_1_q_reg_7_ ( .D(n2453), .CK(CLK), .RN(RST_n), .Q(mul1_reg[7]), 
        .QN(n2192) );
  DFFR_X1 REG1_1_q_reg_8_ ( .D(n2452), .CK(CLK), .RN(RST_n), .Q(mul1_reg[8]), 
        .QN(n2191) );
  DFFR_X1 REG1_1_q_reg_9_ ( .D(n2451), .CK(CLK), .RN(RST_n), .Q(mul1_reg[9]), 
        .QN(n2190) );
  DFFR_X1 REG1_1_q_reg_10_ ( .D(n2450), .CK(CLK), .RN(RST_n), .Q(mul1_reg[10]), 
        .QN(n2189) );
  DFFR_X1 REG1_1_q_reg_11_ ( .D(n2449), .CK(CLK), .RN(RST_n), .Q(mul1_reg[11]), 
        .QN(n2188) );
  DFFR_X1 REG1_1_q_reg_12_ ( .D(n2448), .CK(CLK), .RN(RST_n), .Q(mul1_reg[12]), 
        .QN(n2187) );
  DFFR_X1 REG1_1_q_reg_13_ ( .D(n2447), .CK(CLK), .RN(RST_n), .Q(mul1_reg[13]), 
        .QN(n2186) );
  DFFR_X1 REG11_q_reg_13_ ( .D(n2446), .CK(CLK), .RN(RST_n), .Q(reg2[13]), 
        .QN(n2860) );
  DFFR_X1 REGISTER2_q_reg_13_ ( .D(n2445), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[13]), .QN(n2866) );
  DFFR_X1 REG2_1_q_reg_0_ ( .D(n2444), .CK(CLK), .RN(RST_n), .Q(mul2_reg[0]), 
        .QN(n2185) );
  DFFR_X1 REG2_1_q_reg_1_ ( .D(n2443), .CK(CLK), .RN(RST_n), .Q(mul2_reg[1]), 
        .QN(n2184) );
  DFFR_X1 REG2_1_q_reg_2_ ( .D(n2442), .CK(CLK), .RN(RST_n), .Q(mul2_reg[2]), 
        .QN(n2183) );
  DFFR_X1 REG2_1_q_reg_3_ ( .D(n2441), .CK(CLK), .RN(RST_n), .Q(mul2_reg[3]), 
        .QN(n2182) );
  DFFR_X1 REG2_1_q_reg_4_ ( .D(n2440), .CK(CLK), .RN(RST_n), .Q(mul2_reg[4]), 
        .QN(n2181) );
  DFFR_X1 REG2_1_q_reg_5_ ( .D(n2439), .CK(CLK), .RN(RST_n), .Q(mul2_reg[5]), 
        .QN(n2180) );
  DFFR_X1 REG2_1_q_reg_6_ ( .D(n2438), .CK(CLK), .RN(RST_n), .Q(mul2_reg[6]), 
        .QN(n2179) );
  DFFR_X1 REG2_1_q_reg_7_ ( .D(n2437), .CK(CLK), .RN(RST_n), .Q(mul2_reg[7]), 
        .QN(n2178) );
  DFFR_X1 REG2_1_q_reg_8_ ( .D(n2436), .CK(CLK), .RN(RST_n), .Q(mul2_reg[8]), 
        .QN(n2177) );
  DFFR_X1 REG2_1_q_reg_9_ ( .D(n2435), .CK(CLK), .RN(RST_n), .Q(mul2_reg[9]), 
        .QN(n2176) );
  DFFR_X1 REG2_1_q_reg_10_ ( .D(n2434), .CK(CLK), .RN(RST_n), .Q(mul2_reg[10]), 
        .QN(n2175) );
  DFFR_X1 REG2_1_q_reg_11_ ( .D(n2433), .CK(CLK), .RN(RST_n), .Q(mul2_reg[11]), 
        .QN(n2174) );
  DFFR_X1 REG2_1_q_reg_12_ ( .D(n2432), .CK(CLK), .RN(RST_n), .Q(mul2_reg[12]), 
        .QN(n2173) );
  DFFR_X1 REG21_q_reg_13_ ( .D(n2430), .CK(CLK), .RN(RST_n), .QN(n2878) );
  DFFR_X1 REGISTER3_q_reg_13_ ( .D(n2429), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[13]), .QN(n2805) );
  DFFR_X1 REG3_1_q_reg_0_ ( .D(n2428), .CK(CLK), .RN(RST_n), .Q(mul3_reg[0]), 
        .QN(n2170) );
  DFFR_X1 REG3_1_q_reg_1_ ( .D(n2427), .CK(CLK), .RN(RST_n), .Q(mul3_reg[1]), 
        .QN(n2169) );
  DFFR_X1 REG3_1_q_reg_2_ ( .D(n2426), .CK(CLK), .RN(RST_n), .Q(mul3_reg[2]), 
        .QN(n2168) );
  DFFR_X1 REG3_1_q_reg_3_ ( .D(n2425), .CK(CLK), .RN(RST_n), .Q(mul3_reg[3]), 
        .QN(n2167) );
  DFFR_X1 REG3_1_q_reg_4_ ( .D(n2424), .CK(CLK), .RN(RST_n), .Q(mul3_reg[4]), 
        .QN(n2166) );
  DFFR_X1 REG3_1_q_reg_5_ ( .D(n2423), .CK(CLK), .RN(RST_n), .Q(mul3_reg[5]), 
        .QN(n2165) );
  DFFR_X1 REG3_1_q_reg_6_ ( .D(n2422), .CK(CLK), .RN(RST_n), .Q(mul3_reg[6]), 
        .QN(n2164) );
  DFFR_X1 REG3_1_q_reg_7_ ( .D(n2421), .CK(CLK), .RN(RST_n), .Q(mul3_reg[7]), 
        .QN(n2163) );
  DFFR_X1 REG3_1_q_reg_8_ ( .D(n2420), .CK(CLK), .RN(RST_n), .Q(mul3_reg[8]), 
        .QN(n2162) );
  DFFR_X1 REG3_1_q_reg_9_ ( .D(n2419), .CK(CLK), .RN(RST_n), .Q(mul3_reg[9]), 
        .QN(n2161) );
  DFFR_X1 REG3_1_q_reg_10_ ( .D(n2418), .CK(CLK), .RN(RST_n), .Q(mul3_reg[10]), 
        .QN(n2160) );
  DFFR_X1 REG3_1_q_reg_11_ ( .D(n2417), .CK(CLK), .RN(RST_n), .Q(mul3_reg[11]), 
        .QN(n2159) );
  DFFR_X1 REG3_1_q_reg_12_ ( .D(n2416), .CK(CLK), .RN(RST_n), .Q(mul3_reg[12]), 
        .QN(n2158) );
  DFFR_X1 REG31_q_reg_13_ ( .D(n2414), .CK(CLK), .RN(RST_n), .Q(reg4[13]), 
        .QN(n2859) );
  DFFR_X1 REG41_q_reg_13_ ( .D(n2413), .CK(CLK), .RN(RST_n), .QN(n2879) );
  DFFR_X1 REGISTER4_q_reg_13_ ( .D(n2412), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[13]), .QN(n2804) );
  DFFR_X1 REG4_1_q_reg_0_ ( .D(n2411), .CK(CLK), .RN(RST_n), .Q(mul4_reg[0]), 
        .QN(n2155) );
  DFFR_X1 REG4_1_q_reg_1_ ( .D(n2410), .CK(CLK), .RN(RST_n), .Q(mul4_reg[1]), 
        .QN(n2154) );
  DFFR_X1 REG4_1_q_reg_2_ ( .D(n2409), .CK(CLK), .RN(RST_n), .Q(mul4_reg[2]), 
        .QN(n2153) );
  DFFR_X1 REG4_1_q_reg_3_ ( .D(n2408), .CK(CLK), .RN(RST_n), .Q(mul4_reg[3]), 
        .QN(n2152) );
  DFFR_X1 REG4_1_q_reg_4_ ( .D(n2407), .CK(CLK), .RN(RST_n), .Q(mul4_reg[4]), 
        .QN(n2151) );
  DFFR_X1 REG4_1_q_reg_5_ ( .D(n2406), .CK(CLK), .RN(RST_n), .Q(mul4_reg[5]), 
        .QN(n2150) );
  DFFR_X1 REG4_1_q_reg_6_ ( .D(n2405), .CK(CLK), .RN(RST_n), .Q(mul4_reg[6]), 
        .QN(n2149) );
  DFFR_X1 REG4_1_q_reg_7_ ( .D(n2404), .CK(CLK), .RN(RST_n), .Q(mul4_reg[7]), 
        .QN(n2148) );
  DFFR_X1 REG4_1_q_reg_8_ ( .D(n2403), .CK(CLK), .RN(RST_n), .Q(mul4_reg[8]), 
        .QN(n2147) );
  DFFR_X1 REG4_1_q_reg_9_ ( .D(n2402), .CK(CLK), .RN(RST_n), .Q(mul4_reg[9]), 
        .QN(n2146) );
  DFFR_X1 REG4_1_q_reg_10_ ( .D(n2401), .CK(CLK), .RN(RST_n), .Q(mul4_reg[10]), 
        .QN(n2145) );
  DFFR_X1 REG4_1_q_reg_11_ ( .D(n2400), .CK(CLK), .RN(RST_n), .Q(mul4_reg[11]), 
        .QN(n2144) );
  DFFR_X1 REG4_1_q_reg_12_ ( .D(n2399), .CK(CLK), .RN(RST_n), .Q(mul4_reg[12]), 
        .QN(n2143) );
  DFFR_X1 REGISTER_out_q_reg_0_ ( .D(n2397), .CK(CLK), .RN(RST_n), .Q(DOUT[0]), 
        .QN(n2141) );
  DFFR_X1 REGISTER_out_q_reg_1_ ( .D(n2396), .CK(CLK), .RN(RST_n), .Q(DOUT[1]), 
        .QN(n2140) );
  DFFR_X1 REGISTER_out_q_reg_2_ ( .D(n2395), .CK(CLK), .RN(RST_n), .Q(DOUT[2]), 
        .QN(n2139) );
  DFFR_X1 REGISTER_out_q_reg_3_ ( .D(n2394), .CK(CLK), .RN(RST_n), .Q(DOUT[3]), 
        .QN(n2138) );
  DFFR_X1 REGISTER_out_q_reg_4_ ( .D(n2393), .CK(CLK), .RN(RST_n), .Q(DOUT[4]), 
        .QN(n2137) );
  DFFR_X1 REGISTER_out_q_reg_5_ ( .D(n2392), .CK(CLK), .RN(RST_n), .Q(DOUT[5]), 
        .QN(n2136) );
  DFFR_X1 REGISTER_out_q_reg_6_ ( .D(n2391), .CK(CLK), .RN(RST_n), .Q(DOUT[6]), 
        .QN(n2135) );
  DFFR_X1 REGISTER_out_q_reg_7_ ( .D(n2390), .CK(CLK), .RN(RST_n), .Q(DOUT[7]), 
        .QN(n2134) );
  DFFR_X1 REGISTER_out_q_reg_8_ ( .D(n2389), .CK(CLK), .RN(RST_n), .Q(DOUT[8]), 
        .QN(n2133) );
  DFFR_X1 REGISTER_out_q_reg_9_ ( .D(n2388), .CK(CLK), .RN(RST_n), .Q(DOUT[9]), 
        .QN(n2132) );
  DFFR_X1 REGISTER_out_q_reg_10_ ( .D(n2387), .CK(CLK), .RN(RST_n), .Q(
        DOUT[10]), .QN(n2131) );
  DFFR_X1 REGISTER_out_q_reg_11_ ( .D(n2386), .CK(CLK), .RN(RST_n), .Q(
        DOUT[11]), .QN(n2130) );
  DFFR_X1 REGISTER_out_q_reg_12_ ( .D(n2385), .CK(CLK), .RN(RST_n), .Q(
        DOUT[12]), .QN(n2129) );
  DFFR_X1 REGISTER_out_q_reg_13_ ( .D(n2384), .CK(CLK), .RN(RST_n), .Q(
        DOUT[13]), .QN(n2128) );
  DFFR_X1 REG51_q_reg_0_ ( .D(n2383), .CK(CLK), .RN(RST_n), .Q(reg6[0]), .QN(
        n2660) );
  DFFR_X1 REG51_q_reg_1_ ( .D(n2382), .CK(CLK), .RN(RST_n), .Q(reg6[1]), .QN(
        n2672) );
  DFFR_X1 REG51_q_reg_2_ ( .D(n2381), .CK(CLK), .RN(RST_n), .Q(reg6[2]), .QN(
        n2681) );
  DFFR_X1 REG51_q_reg_3_ ( .D(n2380), .CK(CLK), .RN(RST_n), .Q(reg6[3]), .QN(
        n2680) );
  DFFR_X1 REG51_q_reg_4_ ( .D(n2379), .CK(CLK), .RN(RST_n), .Q(reg6[4]), .QN(
        n2679) );
  DFFR_X1 REG51_q_reg_5_ ( .D(n2378), .CK(CLK), .RN(RST_n), .Q(reg6[5]), .QN(
        n2678) );
  DFFR_X1 REG51_q_reg_6_ ( .D(n2377), .CK(CLK), .RN(RST_n), .Q(reg6[6]), .QN(
        n2677) );
  DFFR_X1 REG51_q_reg_7_ ( .D(n2376), .CK(CLK), .RN(RST_n), .Q(reg6[7]), .QN(
        n2676) );
  DFFR_X1 REG51_q_reg_8_ ( .D(n2375), .CK(CLK), .RN(RST_n), .Q(reg6[8]), .QN(
        n2675) );
  DFFR_X1 REG51_q_reg_9_ ( .D(n2374), .CK(CLK), .RN(RST_n), .Q(reg6[9]), .QN(
        n2674) );
  DFFR_X1 REG51_q_reg_10_ ( .D(n2373), .CK(CLK), .RN(RST_n), .Q(reg6[10]), 
        .QN(n2685) );
  DFFR_X1 REG51_q_reg_11_ ( .D(n2372), .CK(CLK), .RN(RST_n), .Q(reg6[11]), 
        .QN(n2684) );
  DFFR_X1 REG51_q_reg_12_ ( .D(n2371), .CK(CLK), .RN(RST_n), .Q(reg6[12]), 
        .QN(n2683) );
  DFFR_X1 REG51_q_reg_13_ ( .D(n2370), .CK(CLK), .RN(RST_n), .Q(reg6[13]) );
  DFFR_X1 REG61_q_reg_0_ ( .D(n2369), .CK(CLK), .RN(RST_n), .Q(reg7[0]), .QN(
        n2673) );
  DFFR_X1 REG61_q_reg_1_ ( .D(n2368), .CK(CLK), .RN(RST_n), .Q(reg7[1]) );
  DFFR_X1 REG61_q_reg_2_ ( .D(n2367), .CK(CLK), .RN(RST_n), .Q(reg7[2]), .QN(
        n2668) );
  DFFR_X1 REG61_q_reg_3_ ( .D(n2366), .CK(CLK), .RN(RST_n), .Q(reg7[3]), .QN(
        n2667) );
  DFFR_X1 REG61_q_reg_4_ ( .D(n2365), .CK(CLK), .RN(RST_n), .Q(reg7[4]), .QN(
        n2666) );
  DFFR_X1 REG61_q_reg_5_ ( .D(n2364), .CK(CLK), .RN(RST_n), .Q(reg7[5]), .QN(
        n2665) );
  DFFR_X1 REG61_q_reg_6_ ( .D(n2363), .CK(CLK), .RN(RST_n), .Q(reg7[6]), .QN(
        n2664) );
  DFFR_X1 REG61_q_reg_7_ ( .D(n2362), .CK(CLK), .RN(RST_n), .Q(reg7[7]), .QN(
        n2663) );
  DFFR_X1 REG61_q_reg_8_ ( .D(n2361), .CK(CLK), .RN(RST_n), .Q(reg7[8]), .QN(
        n2662) );
  DFFR_X1 REG61_q_reg_9_ ( .D(n2360), .CK(CLK), .RN(RST_n), .Q(reg7[9]), .QN(
        n2661) );
  DFFR_X1 REG61_q_reg_10_ ( .D(n2359), .CK(CLK), .RN(RST_n), .Q(reg7[10]), 
        .QN(n2671) );
  DFFR_X1 REG61_q_reg_11_ ( .D(n2358), .CK(CLK), .RN(RST_n), .Q(reg7[11]), 
        .QN(n2670) );
  DFFR_X1 REG61_q_reg_12_ ( .D(n2357), .CK(CLK), .RN(RST_n), .Q(reg7[12]), 
        .QN(n2669) );
  XOR2_X1 U27 ( .A(n23), .B(n24), .Z(n22) );
  XOR2_X1 U32 ( .A(n33), .B(n34), .Z(n32) );
  XOR2_X1 U35 ( .A(n40), .B(n41), .Z(p9_S[67]) );
  XOR2_X1 U38 ( .A(n46), .B(n47), .Z(n45) );
  XOR2_X1 U40 ( .A(n50), .B(n51), .Z(n49) );
  XOR2_X1 U42 ( .A(n54), .B(n55), .Z(n52) );
  XOR2_X1 U44 ( .A(n58), .B(n59), .Z(n57) );
  XOR2_X1 U52 ( .A(n62), .B(n63), .Z(n61) );
  XOR2_X1 U54 ( .A(n66), .B(n67), .Z(n65) );
  XOR2_X1 U56 ( .A(n70), .B(n71), .Z(n69) );
  XOR2_X1 U58 ( .A(n74), .B(n75), .Z(n73) );
  XOR2_X1 U62 ( .A(n82), .B(n83), .Z(n81) );
  XOR2_X1 U92 ( .A(n27), .B(n115), .Z(n118) );
  XOR2_X1 U109 ( .A(n126), .B(n127), .Z(n132) );
  XOR2_X1 U112 ( .A(n137), .B(n123), .Z(n126) );
  XOR2_X1 U125 ( .A(n145), .B(n133), .Z(n129) );
  XOR2_X1 U139 ( .A(n141), .B(n142), .Z(n155) );
  XOR2_X1 U149 ( .A(p9_muxs_out_3__18_), .B(n148), .Z(n161) );
  XOR2_X1 U157 ( .A(n164), .B(n163), .Z(n166) );
  XOR2_X1 U166 ( .A(n157), .B(n175), .Z(n164) );
  XOR2_X1 U167 ( .A(p9_muxs_out_2__17_), .B(p9_muxs_out_3__17_), .Z(n175) );
  XOR2_X1 U173 ( .A(n182), .B(n179), .Z(n55) );
  XOR2_X1 U197 ( .A(n207), .B(n195), .Z(n58) );
  XOR2_X1 U209 ( .A(n187), .B(n188), .Z(n215) );
  XOR2_X1 U221 ( .A(n205), .B(n204), .Z(n227) );
  XOR2_X1 U222 ( .A(n231), .B(n208), .Z(n204) );
  XOR2_X1 U224 ( .A(n232), .B(n218), .Z(n210) );
  XOR2_X1 U228 ( .A(p9_muxs_out_1__14_), .B(n217), .Z(n209) );
  XOR2_X1 U245 ( .A(n225), .B(n224), .Z(n244) );
  XOR2_X1 U246 ( .A(n248), .B(n230), .Z(n224) );
  XOR2_X1 U254 ( .A(p9_muxs_out_3__13_), .B(n238), .Z(n253) );
  XOR2_X1 U273 ( .A(n241), .B(n242), .Z(n265) );
  XOR2_X1 U274 ( .A(n266), .B(n247), .Z(n242) );
  XOR2_X1 U281 ( .A(p9_muxs_out_3__12_), .B(n261), .Z(n270) );
  XOR2_X1 U285 ( .A(n239), .B(n272), .Z(n241) );
  XOR2_X1 U297 ( .A(n262), .B(n263), .Z(n287) );
  XOR2_X1 U321 ( .A(n284), .B(n285), .Z(n301) );
  XOR2_X1 U330 ( .A(n282), .B(n283), .Z(n284) );
  XOR2_X1 U344 ( .A(p9_muxs_out_3__9_), .B(n300), .Z(n310) );
  XOR2_X1 U361 ( .A(n322), .B(n323), .Z(n327) );
  XOR2_X1 U362 ( .A(p9_muxs_out_3__8_), .B(n321), .Z(n322) );
  XOR2_X1 U380 ( .A(p9_muxs_out_2__7_), .B(n325), .Z(n331) );
  XOR2_X1 U409 ( .A(n349), .B(n350), .Z(n348) );
  XOR2_X1 U414 ( .A(n359), .B(n360), .Z(n358) );
  XOR2_X1 U417 ( .A(n366), .B(n367), .Z(p8_S[67]) );
  XOR2_X1 U420 ( .A(n372), .B(n373), .Z(n371) );
  XOR2_X1 U422 ( .A(n376), .B(n377), .Z(n375) );
  XOR2_X1 U424 ( .A(n380), .B(n381), .Z(n378) );
  XOR2_X1 U426 ( .A(n384), .B(n385), .Z(n383) );
  XOR2_X1 U428 ( .A(n388), .B(n389), .Z(n387) );
  XOR2_X1 U430 ( .A(n392), .B(n393), .Z(n391) );
  XOR2_X1 U432 ( .A(n396), .B(n397), .Z(n395) );
  XOR2_X1 U434 ( .A(n400), .B(n401), .Z(n399) );
  XOR2_X1 U438 ( .A(n408), .B(n409), .Z(n407) );
  XOR2_X1 U468 ( .A(n353), .B(n441), .Z(n444) );
  XOR2_X1 U485 ( .A(n452), .B(n453), .Z(n458) );
  XOR2_X1 U488 ( .A(n463), .B(n449), .Z(n452) );
  XOR2_X1 U501 ( .A(n471), .B(n459), .Z(n455) );
  XOR2_X1 U515 ( .A(n467), .B(n468), .Z(n481) );
  XOR2_X1 U525 ( .A(p8_muxs_out_3__18_), .B(n474), .Z(n487) );
  XOR2_X1 U533 ( .A(n490), .B(n489), .Z(n492) );
  XOR2_X1 U542 ( .A(n483), .B(n501), .Z(n490) );
  XOR2_X1 U543 ( .A(p8_muxs_out_2__17_), .B(p8_muxs_out_3__17_), .Z(n501) );
  XOR2_X1 U549 ( .A(n508), .B(n505), .Z(n381) );
  XOR2_X1 U573 ( .A(n533), .B(n521), .Z(n384) );
  XOR2_X1 U585 ( .A(n513), .B(n514), .Z(n541) );
  XOR2_X1 U597 ( .A(n531), .B(n530), .Z(n553) );
  XOR2_X1 U598 ( .A(n557), .B(n534), .Z(n530) );
  XOR2_X1 U600 ( .A(n558), .B(n544), .Z(n536) );
  XOR2_X1 U604 ( .A(p8_muxs_out_1__14_), .B(n543), .Z(n535) );
  XOR2_X1 U621 ( .A(n551), .B(n550), .Z(n570) );
  XOR2_X1 U622 ( .A(n574), .B(n556), .Z(n550) );
  XOR2_X1 U630 ( .A(p8_muxs_out_3__13_), .B(n564), .Z(n579) );
  XOR2_X1 U649 ( .A(n567), .B(n568), .Z(n591) );
  XOR2_X1 U650 ( .A(n592), .B(n573), .Z(n568) );
  XOR2_X1 U657 ( .A(p8_muxs_out_3__12_), .B(n587), .Z(n596) );
  XOR2_X1 U661 ( .A(n565), .B(n598), .Z(n567) );
  XOR2_X1 U673 ( .A(n588), .B(n589), .Z(n613) );
  XOR2_X1 U697 ( .A(n610), .B(n611), .Z(n627) );
  XOR2_X1 U706 ( .A(n608), .B(n609), .Z(n610) );
  XOR2_X1 U720 ( .A(p8_muxs_out_3__9_), .B(n626), .Z(n636) );
  XOR2_X1 U737 ( .A(n648), .B(n649), .Z(n653) );
  XOR2_X1 U738 ( .A(p8_muxs_out_3__8_), .B(n647), .Z(n648) );
  XOR2_X1 U756 ( .A(p8_muxs_out_2__7_), .B(n651), .Z(n657) );
  XOR2_X1 U785 ( .A(n675), .B(n676), .Z(n674) );
  XOR2_X1 U790 ( .A(n685), .B(n686), .Z(n684) );
  XOR2_X1 U793 ( .A(n692), .B(n693), .Z(p7_S[67]) );
  XOR2_X1 U796 ( .A(n698), .B(n699), .Z(n697) );
  XOR2_X1 U798 ( .A(n702), .B(n703), .Z(n701) );
  XOR2_X1 U800 ( .A(n706), .B(n707), .Z(n704) );
  XOR2_X1 U802 ( .A(n710), .B(n711), .Z(n709) );
  XOR2_X1 U804 ( .A(n714), .B(n715), .Z(n713) );
  XOR2_X1 U806 ( .A(n718), .B(n719), .Z(n717) );
  XOR2_X1 U808 ( .A(n722), .B(n723), .Z(n721) );
  XOR2_X1 U810 ( .A(n726), .B(n727), .Z(n725) );
  XOR2_X1 U814 ( .A(n734), .B(n735), .Z(n733) );
  XOR2_X1 U844 ( .A(n679), .B(n767), .Z(n770) );
  XOR2_X1 U861 ( .A(n778), .B(n779), .Z(n784) );
  XOR2_X1 U864 ( .A(n789), .B(n775), .Z(n778) );
  XOR2_X1 U877 ( .A(n797), .B(n785), .Z(n781) );
  XOR2_X1 U891 ( .A(n793), .B(n794), .Z(n807) );
  XOR2_X1 U901 ( .A(p7_muxs_out_3__18_), .B(n800), .Z(n813) );
  XOR2_X1 U909 ( .A(n816), .B(n815), .Z(n818) );
  XOR2_X1 U918 ( .A(n809), .B(n827), .Z(n816) );
  XOR2_X1 U919 ( .A(p7_muxs_out_2__17_), .B(p7_muxs_out_3__17_), .Z(n827) );
  XOR2_X1 U925 ( .A(n834), .B(n831), .Z(n707) );
  XOR2_X1 U949 ( .A(n859), .B(n847), .Z(n710) );
  XOR2_X1 U961 ( .A(n839), .B(n840), .Z(n867) );
  XOR2_X1 U973 ( .A(n857), .B(n856), .Z(n879) );
  XOR2_X1 U974 ( .A(n883), .B(n860), .Z(n856) );
  XOR2_X1 U976 ( .A(n884), .B(n870), .Z(n862) );
  XOR2_X1 U980 ( .A(p7_muxs_out_1__14_), .B(n869), .Z(n861) );
  XOR2_X1 U997 ( .A(n877), .B(n876), .Z(n896) );
  XOR2_X1 U998 ( .A(n900), .B(n882), .Z(n876) );
  XOR2_X1 U1006 ( .A(p7_muxs_out_3__13_), .B(n890), .Z(n905) );
  XOR2_X1 U1025 ( .A(n893), .B(n894), .Z(n917) );
  XOR2_X1 U1026 ( .A(n918), .B(n899), .Z(n894) );
  XOR2_X1 U1033 ( .A(p7_muxs_out_3__12_), .B(n913), .Z(n922) );
  XOR2_X1 U1037 ( .A(n891), .B(n924), .Z(n893) );
  XOR2_X1 U1049 ( .A(n914), .B(n915), .Z(n939) );
  XOR2_X1 U1073 ( .A(n936), .B(n937), .Z(n953) );
  XOR2_X1 U1082 ( .A(n934), .B(n935), .Z(n936) );
  XOR2_X1 U1096 ( .A(p7_muxs_out_3__9_), .B(n952), .Z(n962) );
  XOR2_X1 U1113 ( .A(n974), .B(n975), .Z(n979) );
  XOR2_X1 U1114 ( .A(p7_muxs_out_3__8_), .B(n973), .Z(n974) );
  XOR2_X1 U1132 ( .A(p7_muxs_out_2__7_), .B(n977), .Z(n983) );
  XOR2_X1 U1161 ( .A(n1001), .B(n1002), .Z(n1000) );
  XOR2_X1 U1166 ( .A(n1011), .B(n1012), .Z(n1010) );
  XOR2_X1 U1169 ( .A(n1018), .B(n1019), .Z(p6_S[67]) );
  XOR2_X1 U1172 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR2_X1 U1174 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR2_X1 U1176 ( .A(n1032), .B(n1033), .Z(n1030) );
  XOR2_X1 U1178 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR2_X1 U1180 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR2_X1 U1182 ( .A(n1044), .B(n1045), .Z(n1043) );
  XOR2_X1 U1184 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR2_X1 U1186 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR2_X1 U1188 ( .A(n1056), .B(n1057), .Z(n1055) );
  XOR2_X1 U1190 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR2_X1 U1220 ( .A(n1005), .B(n1093), .Z(n1096) );
  XOR2_X1 U1237 ( .A(n1104), .B(n1105), .Z(n1110) );
  XOR2_X1 U1240 ( .A(n1115), .B(n1101), .Z(n1104) );
  XOR2_X1 U1253 ( .A(n1123), .B(n1111), .Z(n1107) );
  XOR2_X1 U1267 ( .A(n1119), .B(n1120), .Z(n1133) );
  XOR2_X1 U1277 ( .A(p6_muxs_out_3__18_), .B(n1126), .Z(n1139) );
  XOR2_X1 U1285 ( .A(n1142), .B(n1141), .Z(n1144) );
  XOR2_X1 U1294 ( .A(n1135), .B(n1153), .Z(n1142) );
  XOR2_X1 U1295 ( .A(p6_muxs_out_2__17_), .B(p6_muxs_out_3__17_), .Z(n1153) );
  XOR2_X1 U1301 ( .A(n1160), .B(n1157), .Z(n1033) );
  XOR2_X1 U1325 ( .A(n1185), .B(n1173), .Z(n1036) );
  XOR2_X1 U1337 ( .A(n1165), .B(n1166), .Z(n1193) );
  XOR2_X1 U1349 ( .A(n1183), .B(n1182), .Z(n1205) );
  XOR2_X1 U1350 ( .A(n1209), .B(n1186), .Z(n1182) );
  XOR2_X1 U1352 ( .A(n1210), .B(n1196), .Z(n1188) );
  XOR2_X1 U1356 ( .A(p6_muxs_out_1__14_), .B(n1195), .Z(n1187) );
  XOR2_X1 U1373 ( .A(n1203), .B(n1202), .Z(n1222) );
  XOR2_X1 U1374 ( .A(n1226), .B(n1208), .Z(n1202) );
  XOR2_X1 U1382 ( .A(p6_muxs_out_3__13_), .B(n1216), .Z(n1231) );
  XOR2_X1 U1401 ( .A(n1219), .B(n1220), .Z(n1243) );
  XOR2_X1 U1402 ( .A(n1244), .B(n1225), .Z(n1220) );
  XOR2_X1 U1409 ( .A(p6_muxs_out_3__12_), .B(n1239), .Z(n1248) );
  XOR2_X1 U1413 ( .A(n1217), .B(n1250), .Z(n1219) );
  XOR2_X1 U1425 ( .A(n1240), .B(n1241), .Z(n1265) );
  XOR2_X1 U1449 ( .A(n1262), .B(n1263), .Z(n1279) );
  XOR2_X1 U1458 ( .A(n1260), .B(n1261), .Z(n1262) );
  XOR2_X1 U1472 ( .A(p6_muxs_out_3__9_), .B(n1278), .Z(n1288) );
  XOR2_X1 U1489 ( .A(n1300), .B(n1301), .Z(n1305) );
  XOR2_X1 U1490 ( .A(p6_muxs_out_3__8_), .B(n1299), .Z(n1300) );
  XOR2_X1 U1508 ( .A(p6_muxs_out_2__7_), .B(n1303), .Z(n1309) );
  XOR2_X1 U1537 ( .A(n1329), .B(n1330), .Z(n1328) );
  XOR2_X1 U1542 ( .A(n1339), .B(n1340), .Z(n1338) );
  XOR2_X1 U1545 ( .A(n1346), .B(n1347), .Z(p11_S[67]) );
  XOR2_X1 U1548 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR2_X1 U1550 ( .A(n1356), .B(n1357), .Z(n1355) );
  XOR2_X1 U1552 ( .A(n1360), .B(n1361), .Z(n1358) );
  XOR2_X1 U1554 ( .A(n1364), .B(n1365), .Z(n1363) );
  XOR2_X1 U1556 ( .A(n1368), .B(n1369), .Z(n1367) );
  XOR2_X1 U1558 ( .A(n1372), .B(n1373), .Z(n1371) );
  XOR2_X1 U1560 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR2_X1 U1562 ( .A(n1380), .B(n1381), .Z(n1379) );
  XOR2_X1 U1566 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR2_X1 U1596 ( .A(n1333), .B(n1424), .Z(n1427) );
  XOR2_X1 U1613 ( .A(n1436), .B(n1437), .Z(n1442) );
  XOR2_X1 U1616 ( .A(n1448), .B(n1432), .Z(n1436) );
  XOR2_X1 U1627 ( .A(n1457), .B(n1443), .Z(n1439) );
  XOR2_X1 U1640 ( .A(n1453), .B(n1454), .Z(n1467) );
  XOR2_X1 U1650 ( .A(p11_muxs_out_3__18_), .B(n1460), .Z(n1474) );
  XOR2_X1 U1658 ( .A(n1477), .B(n1476), .Z(n1479) );
  XOR2_X1 U1667 ( .A(n1469), .B(n1489), .Z(n1477) );
  XOR2_X1 U1668 ( .A(p11_muxs_out_2__17_), .B(p11_muxs_out_3__17_), .Z(n1489)
         );
  XOR2_X1 U1674 ( .A(n1496), .B(n1493), .Z(n1361) );
  XOR2_X1 U1698 ( .A(n1522), .B(n1510), .Z(n1364) );
  XOR2_X1 U1710 ( .A(n1501), .B(n1502), .Z(n1531) );
  XOR2_X1 U1721 ( .A(n1520), .B(n1519), .Z(n1542) );
  XOR2_X1 U1722 ( .A(n1546), .B(n1523), .Z(n1519) );
  XOR2_X1 U1724 ( .A(n1547), .B(n1534), .Z(n1525) );
  XOR2_X1 U1728 ( .A(p11_muxs_out_1__14_), .B(n1533), .Z(n1524) );
  XOR2_X1 U1745 ( .A(n1540), .B(n1539), .Z(n1561) );
  XOR2_X1 U1747 ( .A(n1544), .B(n1545), .Z(n1565) );
  XOR2_X1 U1752 ( .A(p11_muxs_out_2__13_), .B(n1570), .Z(n1543) );
  XOR2_X1 U1757 ( .A(n1537), .B(n1535), .Z(n1572) );
  XOR2_X1 U1777 ( .A(p11_muxs_out_3__12_), .B(n1580), .Z(n1586) );
  XOR2_X1 U1785 ( .A(n1555), .B(n1592), .Z(n1558) );
  XOR2_X1 U1798 ( .A(n1581), .B(n1582), .Z(n1605) );
  XOR2_X1 U1829 ( .A(n1600), .B(n1601), .Z(n1602) );
  XOR2_X1 U1842 ( .A(p11_muxs_out_3__9_), .B(n1617), .Z(n1627) );
  XOR2_X1 U1857 ( .A(n1639), .B(n1640), .Z(n1644) );
  XOR2_X1 U1858 ( .A(p11_muxs_out_3__8_), .B(n1638), .Z(n1639) );
  XOR2_X1 U1875 ( .A(p11_muxs_out_2__7_), .B(n1642), .Z(n1648) );
  XOR2_X1 U1904 ( .A(n1669), .B(n1670), .Z(n1668) );
  XOR2_X1 U1909 ( .A(n1679), .B(n1680), .Z(n1678) );
  XOR2_X1 U1912 ( .A(n1686), .B(n1687), .Z(p10_S[67]) );
  XOR2_X1 U1915 ( .A(n1692), .B(n1693), .Z(n1691) );
  XOR2_X1 U1917 ( .A(n1696), .B(n1697), .Z(n1695) );
  XOR2_X1 U1919 ( .A(n1700), .B(n1701), .Z(n1698) );
  XOR2_X1 U1921 ( .A(n1704), .B(n1705), .Z(n1703) );
  XOR2_X1 U1923 ( .A(n1708), .B(n1709), .Z(n1707) );
  XOR2_X1 U1925 ( .A(n1712), .B(n1713), .Z(n1711) );
  XOR2_X1 U1927 ( .A(n1716), .B(n1717), .Z(n1715) );
  XOR2_X1 U1929 ( .A(n1720), .B(n1721), .Z(n1719) );
  XOR2_X1 U1933 ( .A(n1728), .B(n1729), .Z(n1727) );
  XOR2_X1 U1963 ( .A(n1673), .B(n1764), .Z(n1767) );
  XOR2_X1 U1980 ( .A(n1776), .B(n1777), .Z(n1782) );
  XOR2_X1 U1983 ( .A(n1788), .B(n1772), .Z(n1776) );
  XOR2_X1 U1994 ( .A(n1797), .B(n1783), .Z(n1779) );
  XOR2_X1 U2007 ( .A(n1793), .B(n1794), .Z(n1807) );
  XOR2_X1 U2017 ( .A(p10_muxs_out_3__18_), .B(n1800), .Z(n1814) );
  XOR2_X1 U2025 ( .A(n1817), .B(n1816), .Z(n1819) );
  XOR2_X1 U2034 ( .A(n1809), .B(n1829), .Z(n1817) );
  XOR2_X1 U2035 ( .A(p10_muxs_out_2__17_), .B(p10_muxs_out_3__17_), .Z(n1829)
         );
  XOR2_X1 U2041 ( .A(n1836), .B(n1833), .Z(n1701) );
  XOR2_X1 U2065 ( .A(n1862), .B(n1850), .Z(n1704) );
  XOR2_X1 U2077 ( .A(n1841), .B(n1842), .Z(n1871) );
  XOR2_X1 U2088 ( .A(n1860), .B(n1859), .Z(n1882) );
  XOR2_X1 U2089 ( .A(n1886), .B(n1863), .Z(n1859) );
  XOR2_X1 U2091 ( .A(n1887), .B(n1874), .Z(n1865) );
  XOR2_X1 U2095 ( .A(p10_muxs_out_1__14_), .B(n1873), .Z(n1864) );
  XOR2_X1 U2112 ( .A(n1880), .B(n1879), .Z(n1901) );
  XOR2_X1 U2114 ( .A(n1884), .B(n1885), .Z(n1905) );
  XOR2_X1 U2119 ( .A(p10_muxs_out_2__13_), .B(n1910), .Z(n1883) );
  XOR2_X1 U2124 ( .A(n1877), .B(n1875), .Z(n1912) );
  XOR2_X1 U2141 ( .A(n1898), .B(n1899), .Z(n1924) );
  XOR2_X1 U2144 ( .A(p10_muxs_out_3__12_), .B(n1920), .Z(n1926) );
  XOR2_X1 U2152 ( .A(n1895), .B(n1932), .Z(n1898) );
  XOR2_X1 U2165 ( .A(n1921), .B(n1922), .Z(n1945) );
  XOR2_X1 U2196 ( .A(n1940), .B(n1941), .Z(n1942) );
  XOR2_X1 U2209 ( .A(p10_muxs_out_3__9_), .B(n1957), .Z(n1967) );
  XOR2_X1 U2224 ( .A(n1979), .B(n1980), .Z(n1984) );
  XOR2_X1 U2225 ( .A(p10_muxs_out_3__8_), .B(n1978), .Z(n1979) );
  XOR2_X1 U2242 ( .A(p10_muxs_out_2__7_), .B(n1982), .Z(n1988) );
  MUX2_X1 U2264 ( .A(reg7[12]), .B(temp6[12]), .S(VIN), .Z(n2357) );
  MUX2_X1 U2265 ( .A(reg7[11]), .B(temp6[11]), .S(VIN), .Z(n2358) );
  MUX2_X1 U2266 ( .A(reg7[10]), .B(temp6[10]), .S(VIN), .Z(n2359) );
  MUX2_X1 U2267 ( .A(reg7[9]), .B(temp6[9]), .S(VIN), .Z(n2360) );
  MUX2_X1 U2268 ( .A(reg7[8]), .B(temp6[8]), .S(VIN), .Z(n2361) );
  MUX2_X1 U2269 ( .A(reg7[7]), .B(temp6[7]), .S(VIN), .Z(n2362) );
  MUX2_X1 U2270 ( .A(reg7[6]), .B(temp6[6]), .S(VIN), .Z(n2363) );
  MUX2_X1 U2271 ( .A(reg7[5]), .B(temp6[5]), .S(VIN), .Z(n2364) );
  MUX2_X1 U2272 ( .A(reg7[4]), .B(temp6[4]), .S(VIN), .Z(n2365) );
  MUX2_X1 U2273 ( .A(reg7[3]), .B(temp6[3]), .S(VIN), .Z(n2366) );
  MUX2_X1 U2274 ( .A(reg7[2]), .B(temp6[2]), .S(VIN), .Z(n2367) );
  MUX2_X1 U2275 ( .A(reg7[1]), .B(temp6[1]), .S(VIN), .Z(n2368) );
  MUX2_X1 U2276 ( .A(reg7[0]), .B(temp6[0]), .S(VIN), .Z(n2369) );
  MUX2_X1 U2277 ( .A(reg6[13]), .B(temp5[13]), .S(VIN), .Z(n2370) );
  MUX2_X1 U2278 ( .A(reg6[12]), .B(temp5[12]), .S(VIN), .Z(n2371) );
  MUX2_X1 U2279 ( .A(reg6[11]), .B(temp5[11]), .S(VIN), .Z(n2372) );
  MUX2_X1 U2280 ( .A(reg6[10]), .B(temp5[10]), .S(VIN), .Z(n2373) );
  MUX2_X1 U2281 ( .A(reg6[9]), .B(temp5[9]), .S(VIN), .Z(n2374) );
  MUX2_X1 U2282 ( .A(reg6[8]), .B(temp5[8]), .S(VIN), .Z(n2375) );
  MUX2_X1 U2283 ( .A(reg6[7]), .B(temp5[7]), .S(VIN), .Z(n2376) );
  MUX2_X1 U2284 ( .A(reg6[6]), .B(temp5[6]), .S(VIN), .Z(n2377) );
  MUX2_X1 U2285 ( .A(reg6[5]), .B(temp5[5]), .S(VIN), .Z(n2378) );
  MUX2_X1 U2286 ( .A(reg6[4]), .B(temp5[4]), .S(VIN), .Z(n2379) );
  MUX2_X1 U2287 ( .A(reg6[3]), .B(temp5[3]), .S(VIN), .Z(n2380) );
  MUX2_X1 U2288 ( .A(reg6[2]), .B(temp5[2]), .S(VIN), .Z(n2381) );
  MUX2_X1 U2289 ( .A(reg6[1]), .B(temp5[1]), .S(VIN), .Z(n2382) );
  MUX2_X1 U2290 ( .A(reg6[0]), .B(temp5[0]), .S(VIN), .Z(n2383) );
  MUX2_X1 U2550 ( .A(reg4_reg[6]), .B(n2212), .S(VIN), .Z(n2510) );
  MUX2_X1 U2555 ( .A(reg3_reg[6]), .B(n2213), .S(VIN), .Z(n2513) );
  MUX2_X1 U2558 ( .A(reg2_reg[6]), .B(reg2[6]), .S(VIN), .Z(n2515) );
  MUX2_X1 U2562 ( .A(reg1_reg[6]), .B(w[6]), .S(VIN), .Z(n2517) );
  MUX2_X1 U2563 ( .A(reg4_reg[5]), .B(n2214), .S(VIN), .Z(n2518) );
  MUX2_X1 U2568 ( .A(reg3_reg[5]), .B(n2215), .S(VIN), .Z(n2521) );
  MUX2_X1 U2571 ( .A(reg2_reg[5]), .B(reg2[5]), .S(VIN), .Z(n2523) );
  MUX2_X1 U2575 ( .A(reg1_reg[5]), .B(w[5]), .S(VIN), .Z(n2525) );
  MUX2_X1 U2588 ( .A(reg1_reg[4]), .B(w[4]), .S(VIN), .Z(n2533) );
  MUX2_X1 U2589 ( .A(reg4_reg[3]), .B(n2218), .S(VIN), .Z(n2534) );
  MUX2_X1 U2594 ( .A(reg3_reg[3]), .B(n2219), .S(VIN), .Z(n2537) );
  MUX2_X1 U2597 ( .A(reg2_reg[3]), .B(reg2[3]), .S(VIN), .Z(n2539) );
  MUX2_X1 U2601 ( .A(reg1_reg[3]), .B(w[3]), .S(VIN), .Z(n2541) );
  MUX2_X1 U2602 ( .A(reg4_reg[2]), .B(n2220), .S(VIN), .Z(n2542) );
  MUX2_X1 U2607 ( .A(reg3_reg[2]), .B(n2221), .S(VIN), .Z(n2545) );
  MUX2_X1 U2610 ( .A(reg2_reg[2]), .B(reg2[2]), .S(VIN), .Z(n2547) );
  MUX2_X1 U2614 ( .A(reg1_reg[2]), .B(w[2]), .S(VIN), .Z(n2549) );
  MUX2_X1 U2651 ( .A(xin[13]), .B(n2240), .S(VIN), .Z(n2567) );
  MUX2_X1 U2652 ( .A(xin[12]), .B(n2239), .S(VIN), .Z(n2568) );
  MUX2_X1 U2653 ( .A(xin[11]), .B(n2238), .S(VIN), .Z(n2569) );
  MUX2_X1 U2654 ( .A(xin[10]), .B(n2237), .S(VIN), .Z(n2570) );
  MUX2_X1 U2655 ( .A(xin[9]), .B(n2236), .S(VIN), .Z(n2571) );
  MUX2_X1 U2656 ( .A(xin[8]), .B(n2235), .S(VIN), .Z(n2572) );
  MUX2_X1 U2657 ( .A(xin[7]), .B(n2234), .S(VIN), .Z(n2573) );
  MUX2_X1 U2658 ( .A(xin[6]), .B(n2233), .S(VIN), .Z(n2574) );
  MUX2_X1 U2659 ( .A(xin[5]), .B(n2232), .S(VIN), .Z(n2575) );
  MUX2_X1 U2660 ( .A(xin[4]), .B(n2231), .S(VIN), .Z(n2576) );
  MUX2_X1 U2661 ( .A(xin[3]), .B(n2230), .S(VIN), .Z(n2577) );
  MUX2_X1 U2662 ( .A(xin[2]), .B(n2229), .S(VIN), .Z(n2578) );
  MUX2_X1 U2663 ( .A(xin[1]), .B(n2228), .S(VIN), .Z(n2579) );
  MUX2_X1 U2664 ( .A(xin[0]), .B(n2227), .S(VIN), .Z(n2580) );
  MUX2_X1 U2667 ( .A(n2227), .B(DIN[0]), .S(VIN), .Z(n2582) );
  MUX2_X1 U2668 ( .A(n2228), .B(DIN[1]), .S(VIN), .Z(n2583) );
  MUX2_X1 U2669 ( .A(n2229), .B(DIN[2]), .S(VIN), .Z(n2584) );
  MUX2_X1 U2670 ( .A(n2230), .B(DIN[3]), .S(VIN), .Z(n2585) );
  MUX2_X1 U2671 ( .A(n2231), .B(DIN[4]), .S(VIN), .Z(n2586) );
  MUX2_X1 U2672 ( .A(n2232), .B(DIN[5]), .S(VIN), .Z(n2587) );
  MUX2_X1 U2673 ( .A(n2233), .B(DIN[6]), .S(VIN), .Z(n2588) );
  MUX2_X1 U2674 ( .A(n2234), .B(DIN[7]), .S(VIN), .Z(n2589) );
  MUX2_X1 U2675 ( .A(n2235), .B(DIN[8]), .S(VIN), .Z(n2590) );
  MUX2_X1 U2676 ( .A(n2236), .B(DIN[9]), .S(VIN), .Z(n2591) );
  MUX2_X1 U2677 ( .A(n2237), .B(DIN[10]), .S(VIN), .Z(n2592) );
  MUX2_X1 U2678 ( .A(n2238), .B(DIN[11]), .S(VIN), .Z(n2593) );
  MUX2_X1 U2679 ( .A(n2239), .B(DIN[12]), .S(VIN), .Z(n2594) );
  MUX2_X1 U2680 ( .A(n2240), .B(DIN[13]), .S(VIN), .Z(n2595) );
  DFFR_X1 REG11_q_reg_12_ ( .D(n2468), .CK(CLK), .RN(RST_n), .Q(reg2[12]), 
        .QN(n2863) );
  DFFR_X1 REG11_q_reg_11_ ( .D(n2476), .CK(CLK), .RN(RST_n), .Q(reg2[11]), 
        .QN(n2862) );
  DFFR_X1 REG31_q_reg_11_ ( .D(n2472), .CK(CLK), .RN(RST_n), .Q(reg4[11]), 
        .QN(n2861) );
  DFFR_X2 REGISTER4_q_reg_5_ ( .D(n2518), .CK(CLK), .RN(RST_n), .Q(reg4_reg[5]), .QN(n2854) );
  DFFR_X2 REGISTER3_q_reg_5_ ( .D(n2521), .CK(CLK), .RN(RST_n), .Q(reg3_reg[5]), .QN(n2853) );
  DFFR_X2 REGISTER2_q_reg_5_ ( .D(n2523), .CK(CLK), .RN(RST_n), .Q(reg2_reg[5]), .QN(n2852) );
  DFFR_X2 REGISTER1_q_reg_5_ ( .D(n2525), .CK(CLK), .RN(RST_n), .Q(reg1_reg[5]), .QN(n2851) );
  DFFR_X2 REGISTER4_q_reg_3_ ( .D(n2534), .CK(CLK), .RN(RST_n), .Q(reg4_reg[3]), .QN(n2847) );
  DFFR_X2 REGISTER3_q_reg_3_ ( .D(n2537), .CK(CLK), .RN(RST_n), .Q(reg3_reg[3]), .QN(n2846) );
  DFFR_X2 REGISTER2_q_reg_3_ ( .D(n2539), .CK(CLK), .RN(RST_n), .Q(reg2_reg[3]), .QN(n2845) );
  DFFR_X2 REGISTER1_q_reg_3_ ( .D(n2541), .CK(CLK), .RN(RST_n), .Q(reg1_reg[3]), .QN(n2844) );
  DFFR_X1 REG11_q_reg_6_ ( .D(n2516), .CK(CLK), .RN(RST_n), .Q(reg2[6]), .QN(
        n2835) );
  DFFR_X1 REG11_q_reg_5_ ( .D(n2524), .CK(CLK), .RN(RST_n), .Q(reg2[5]), .QN(
        n2834) );
  DFFR_X1 REG11_q_reg_10_ ( .D(n2484), .CK(CLK), .RN(RST_n), .Q(reg2[10]), 
        .QN(n2833) );
  DFFR_X1 REG31_q_reg_8_ ( .D(n2496), .CK(CLK), .RN(RST_n), .Q(reg4[8]), .QN(
        n2832) );
  DFFR_X1 REG11_q_reg_7_ ( .D(n2508), .CK(CLK), .RN(RST_n), .Q(reg2[7]), .QN(
        n2831) );
  DFFR_X1 REG31_q_reg_7_ ( .D(n2504), .CK(CLK), .RN(RST_n), .Q(reg4[7]), .QN(
        n2830) );
  DFFR_X1 REG2_1_q_reg_13_ ( .D(n2431), .CK(CLK), .RN(RST_n), .Q(mul2_reg[13]), 
        .QN(n2172) );
  DFFR_X1 REG4_1_q_reg_13_ ( .D(n2398), .CK(CLK), .RN(RST_n), .Q(mul4_reg[13]), 
        .QN(n2142) );
  DFFR_X1 REG3_1_q_reg_13_ ( .D(n2415), .CK(CLK), .RN(RST_n), .Q(mul3_reg[13]), 
        .QN(n2157) );
  DFFR_X1 REGISTER4_q_reg_4_ ( .D(n2526), .CK(CLK), .RN(RST_n), .Q(reg4_reg[4]), .QN(n2829) );
  DFFR_X1 REGISTER3_q_reg_4_ ( .D(n2529), .CK(CLK), .RN(RST_n), .Q(reg3_reg[4]), .QN(n2828) );
  AOI21_X1 U1766 ( .B1(n1578), .B2(n1579), .A(n1326), .ZN(n1576) );
  AOI22_X1 U1787 ( .A1(A1[11]), .A2(n1579), .B1(A1[12]), .B2(n1578), .ZN(n1575) );
  AOI22_X1 U1533 ( .A1(reg2[13]), .A2(n1323), .B1(n1324), .B2(n2860), .ZN(
        n1322) );
  OAI221_X1 U1532 ( .B1(reg2[12]), .B2(n1319), .C1(n2863), .C2(n1321), .A(
        n1322), .ZN(p11_final_product2_26_) );
  AOI22_X1 U1575 ( .A1(reg2[12]), .A2(n1323), .B1(n1324), .B2(n2863), .ZN(
        n1402) );
  OAI221_X1 U1589 ( .B1(reg2[11]), .B2(n1403), .C1(n2862), .C2(n1404), .A(
        n1423), .ZN(n1413) );
  OAI221_X1 U1588 ( .B1(reg2[13]), .B2(n1420), .C1(n2860), .C2(n1421), .A(
        n1422), .ZN(n1416) );
  AOI22_X1 U1586 ( .A1(reg2[10]), .A2(n1323), .B1(n1324), .B2(n2833), .ZN(
        n1419) );
  OAI221_X1 U1585 ( .B1(reg2[9]), .B2(n1319), .C1(n2816), .C2(n1321), .A(n1419), .ZN(n1415) );
  AOI222_X1 U1581 ( .A1(n1413), .A2(n1414), .B1(n1413), .B2(n1415), .C1(n1414), 
        .C2(n1415), .ZN(n1329) );
  AOI22_X1 U1580 ( .A1(reg2[11]), .A2(n1411), .B1(n1412), .B2(n2862), .ZN(
        n1410) );
  AOI221_X1 U1579 ( .B1(reg2[10]), .B2(n1326), .C1(n2833), .C2(n1409), .A(
        n1410), .ZN(n1330) );
  OAI221_X1 U1577 ( .B1(reg2[12]), .B2(n1403), .C1(n2863), .C2(n1404), .A(
        n1405), .ZN(n1327) );
  AOI222_X1 U1576 ( .A1(n1329), .A2(n1330), .B1(n1329), .B2(n1327), .C1(n1330), 
        .C2(n1327), .ZN(p11_C[71]) );
  XNOR2_X1 U1536 ( .A(n1327), .B(n1328), .ZN(p11_S[71]) );
  OAI221_X1 U1599 ( .B1(reg2[12]), .B2(n1420), .C1(n2863), .C2(n1421), .A(
        n1422), .ZN(n1333) );
  OAI221_X1 U1597 ( .B1(reg2[10]), .B2(n1403), .C1(n2833), .C2(n1404), .A(
        n1428), .ZN(n1424) );
  OAI221_X1 U1620 ( .B1(reg2[11]), .B2(n1420), .C1(n2862), .C2(n1421), .A(
        n1450), .ZN(n1431) );
  OAI221_X1 U1617 ( .B1(reg2[9]), .B2(n1403), .C1(n2816), .C2(n1404), .A(n1449), .ZN(n1432) );
  AOI222_X1 U1601 ( .A1(n1431), .A2(n1432), .B1(n1431), .B2(n1433), .C1(n1432), 
        .C2(n1433), .ZN(n1426) );
  AOI222_X1 U1591 ( .A1(n1424), .A2(n1336), .B1(n1424), .B2(n1425), .C1(n1336), 
        .C2(n1425), .ZN(n1332) );
  XNOR2_X1 U1587 ( .A(n1413), .B(n1416), .ZN(n1417) );
  XNOR2_X1 U1584 ( .A(n1417), .B(n1415), .ZN(n1335) );
  AOI222_X1 U1583 ( .A1(n1336), .A2(n1332), .B1(n1336), .B2(n1335), .C1(n1332), 
        .C2(n1335), .ZN(p11_C[70]) );
  AOI22_X1 U1539 ( .A1(n1333), .A2(n1334), .B1(n1335), .B2(n1336), .ZN(n1331)
         );
  XNOR2_X1 U1538 ( .A(n1331), .B(n1332), .ZN(p11_S[70]) );
  XNOR2_X1 U1619 ( .A(p11_muxs_out_3__20_), .B(n1431), .ZN(n1448) );
  AOI22_X1 U1615 ( .A1(reg2[8]), .A2(n1323), .B1(n1324), .B2(n2811), .ZN(n1447) );
  OAI221_X1 U1614 ( .B1(reg2[7]), .B2(n1319), .C1(n2831), .C2(n1321), .A(n1447), .ZN(n1437) );
  AOI22_X1 U1629 ( .A1(reg2[8]), .A2(n1404), .B1(n1403), .B2(n2811), .ZN(n1458) );
  OAI221_X1 U1631 ( .B1(reg2[10]), .B2(n1420), .C1(n2833), .C2(n1421), .A(
        n1459), .ZN(n1445) );
  AOI222_X1 U1611 ( .A1(p11_muxs_out_3__19_), .A2(n1443), .B1(
        p11_muxs_out_3__19_), .B2(n1444), .C1(n1443), .C2(n1444), .ZN(n1438)
         );
  AOI222_X1 U1605 ( .A1(n1436), .A2(n1437), .B1(n1436), .B2(n1438), .C1(n1437), 
        .C2(n1438), .ZN(n1339) );
  AOI22_X1 U1604 ( .A1(reg2[9]), .A2(n1411), .B1(n1412), .B2(n2816), .ZN(n1435) );
  AOI221_X1 U1603 ( .B1(reg2[8]), .B2(n1326), .C1(n2811), .C2(n1409), .A(n1435), .ZN(n1340) );
  XNOR2_X1 U1595 ( .A(n1426), .B(n1427), .ZN(n1337) );
  AOI222_X1 U1594 ( .A1(n1339), .A2(n1340), .B1(n1339), .B2(n1337), .C1(n1340), 
        .C2(n1337), .ZN(p11_C[69]) );
  XNOR2_X1 U1541 ( .A(n1337), .B(n1338), .ZN(p11_S[69]) );
  XNOR2_X1 U1610 ( .A(n1442), .B(n1438), .ZN(n1341) );
  XNOR2_X1 U1630 ( .A(p11_muxs_out_3__19_), .B(n1445), .ZN(n1457) );
  OAI221_X1 U1647 ( .B1(reg2[7]), .B2(n1403), .C1(n2831), .C2(n1404), .A(n1473), .ZN(n1462) );
  AOI22_X1 U1645 ( .A1(reg2[6]), .A2(n1323), .B1(n1324), .B2(n2835), .ZN(n1472) );
  OAI221_X1 U1644 ( .B1(reg2[5]), .B2(n1319), .C1(n2834), .C2(n1321), .A(n1472), .ZN(n1463) );
  AOI222_X1 U1636 ( .A1(p11_muxs_out_2__17_), .A2(n1462), .B1(
        p11_muxs_out_2__17_), .B2(n1463), .C1(n1462), .C2(n1463), .ZN(n1440)
         );
  OAI221_X1 U1651 ( .B1(reg2[9]), .B2(n1420), .C1(n2816), .C2(n1421), .A(n1475), .ZN(n1460) );
  AOI222_X1 U1634 ( .A1(p11_muxs_out_3__18_), .A2(n1460), .B1(
        p11_muxs_out_3__18_), .B2(n1461), .C1(n1460), .C2(n1461), .ZN(n1441)
         );
  OAI222_X1 U1608 ( .A1(n1439), .A2(n1440), .B1(n1439), .B2(n1441), .C1(n1440), 
        .C2(n1441), .ZN(n1343) );
  AOI222_X1 U1606 ( .A1(n1341), .A2(n1345), .B1(n1341), .B2(n1344), .C1(n1345), 
        .C2(n1344), .ZN(p11_C[68]) );
  AOI22_X1 U1544 ( .A1(p11_muxs_out_3__19_), .A2(n1343), .B1(n1344), .B2(n1345), .ZN(n1342) );
  XNOR2_X1 U1543 ( .A(n1341), .B(n1342), .ZN(p11_S[68]) );
  XNOR2_X1 U1633 ( .A(n1440), .B(n1441), .ZN(n1456) );
  XNOR2_X1 U1626 ( .A(n1456), .B(n1439), .ZN(n1346) );
  XNOR2_X1 U1646 ( .A(p11_muxs_out_2__17_), .B(n1462), .ZN(n1470) );
  XNOR2_X1 U1643 ( .A(n1470), .B(n1463), .ZN(n1453) );
  AOI222_X1 U1669 ( .A1(p11_muxs_out_2__16_), .A2(p11_muxs_out_3__16_), .B1(
        p11_muxs_out_2__16_), .B2(n1490), .C1(p11_muxs_out_3__16_), .C2(n1490), 
        .ZN(n1469) );
  AOI222_X1 U1641 ( .A1(p11_muxs_out_2__17_), .A2(n1468), .B1(
        p11_muxs_out_2__17_), .B2(n1469), .C1(n1468), .C2(n1469), .ZN(n1454)
         );
  XNOR2_X1 U1649 ( .A(p11_muxs_out_2__18_), .B(n1474), .ZN(n1455) );
  AOI222_X1 U1625 ( .A1(n1453), .A2(n1454), .B1(n1453), .B2(n1455), .C1(n1454), 
        .C2(n1455), .ZN(n1349) );
  OAI22_X1 U1624 ( .A1(n2831), .A2(n1411), .B1(n1412), .B2(reg2[7]), .ZN(n1452) );
  AOI221_X1 U1623 ( .B1(n2835), .B2(n1409), .C1(reg2[6]), .C2(n1326), .A(n1452), .ZN(n1348) );
  AOI222_X1 U1622 ( .A1(n1346), .A2(n1349), .B1(n1346), .B2(n1348), .C1(n1349), 
        .C2(n1348), .ZN(p11_C[67]) );
  XNOR2_X1 U1546 ( .A(n1348), .B(n1349), .ZN(n1347) );
  OAI221_X1 U1665 ( .B1(reg2[6]), .B2(n1403), .C1(n2835), .C2(n1404), .A(n1488), .ZN(n1464) );
  AOI22_X1 U1664 ( .A1(reg2[5]), .A2(n1323), .B1(n1324), .B2(n2834), .ZN(n1487) );
  OAI221_X1 U1663 ( .B1(reg2[4]), .B2(n1319), .C1(n2817), .C2(n1321), .A(n1487), .ZN(n1465) );
  XNOR2_X1 U1662 ( .A(n1464), .B(n1465), .ZN(n1484) );
  OAI221_X1 U1660 ( .B1(reg2[8]), .B2(n1420), .C1(n2811), .C2(n1421), .A(n1485), .ZN(n1466) );
  XNOR2_X1 U1659 ( .A(n1484), .B(n1466), .ZN(n1476) );
  XNOR2_X1 U1680 ( .A(p11_muxs_out_3__16_), .B(p11_muxs_out_2__16_), .ZN(n1499) );
  XNOR2_X1 U1679 ( .A(n1499), .B(p11_muxs_out_1__16_), .ZN(n1480) );
  AOI222_X1 U1676 ( .A1(p11_muxs_out_3__15_), .A2(p11_muxs_out_2__15_), .B1(
        p11_muxs_out_3__15_), .B2(n1498), .C1(p11_muxs_out_2__15_), .C2(n1498), 
        .ZN(n1481) );
  OAI221_X1 U1681 ( .B1(reg2[7]), .B2(n1420), .C1(n2831), .C2(n1421), .A(n1500), .ZN(n1483) );
  AOI222_X1 U1656 ( .A1(n1480), .A2(n1481), .B1(n1480), .B2(n1482), .C1(n1481), 
        .C2(n1482), .ZN(n1478) );
  AOI222_X1 U1653 ( .A1(n1476), .A2(n1477), .B1(n1476), .B2(n1478), .C1(n1477), 
        .C2(n1478), .ZN(n1352) );
  XNOR2_X1 U1639 ( .A(n1455), .B(n1467), .ZN(n1353) );
  AOI222_X1 U1638 ( .A1(n1464), .A2(n1465), .B1(n1464), .B2(n1466), .C1(n1465), 
        .C2(n1466), .ZN(n1350) );
  AOI222_X1 U1637 ( .A1(n1352), .A2(n1353), .B1(n1352), .B2(n1350), .C1(n1353), 
        .C2(n1350), .ZN(p11_C[66]) );
  XNOR2_X1 U1547 ( .A(n1350), .B(n1351), .ZN(p11_S[66]) );
  OAI221_X1 U1689 ( .B1(reg2[5]), .B2(n1403), .C1(n2834), .C2(n1404), .A(n1507), .ZN(n1494) );
  AOI22_X1 U1687 ( .A1(reg2[4]), .A2(n1323), .B1(n1324), .B2(n2817), .ZN(n1506) );
  OAI221_X1 U1686 ( .B1(reg2[3]), .B2(n1319), .C1(p11_minus_A_shifted_16_), 
        .C2(n1321), .A(n1506), .ZN(n1495) );
  AOI222_X1 U1672 ( .A1(p11_muxs_out_1__15_), .A2(n1494), .B1(
        p11_muxs_out_1__15_), .B2(n1495), .C1(n1494), .C2(n1495), .ZN(n1356)
         );
  XNOR2_X1 U1688 ( .A(p11_muxs_out_1__15_), .B(n1494), .ZN(n1504) );
  XNOR2_X1 U1685 ( .A(n1504), .B(n1495), .ZN(n1491) );
  NOR2_X1 U1713 ( .A1(p11_muxs_out_1__14_), .A2(n1533), .ZN(n1501) );
  XNOR2_X1 U1712 ( .A(p11_muxs_out_1__15_), .B(p11_muxs_out_3__15_), .ZN(n1532) );
  XNOR2_X1 U1711 ( .A(n1532), .B(p11_muxs_out_2__15_), .ZN(n1502) );
  OAI221_X1 U1725 ( .B1(reg2[5]), .B2(n1420), .C1(n2834), .C2(n1421), .A(n1548), .ZN(n1534) );
  AOI222_X1 U1714 ( .A1(p11_muxs_out_3__14_), .A2(p11_muxs_out_2__14_), .B1(
        p11_muxs_out_3__14_), .B2(n1534), .C1(p11_muxs_out_2__14_), .C2(n1534), 
        .ZN(n1503) );
  AOI222_X1 U1684 ( .A1(n1501), .A2(n1502), .B1(n1501), .B2(n1503), .C1(n1502), 
        .C2(n1503), .ZN(n1492) );
  XNOR2_X1 U1678 ( .A(n1483), .B(n1480), .ZN(n1497) );
  XNOR2_X1 U1675 ( .A(n1497), .B(n1481), .ZN(n1493) );
  AOI222_X1 U1671 ( .A1(n1491), .A2(n1492), .B1(n1491), .B2(n1493), .C1(n1492), 
        .C2(n1493), .ZN(n1357) );
  XNOR2_X1 U1655 ( .A(n1479), .B(n1478), .ZN(n1354) );
  AOI222_X1 U1654 ( .A1(n1356), .A2(n1357), .B1(n1356), .B2(n1354), .C1(n1357), 
        .C2(n1354), .ZN(p11_C[65]) );
  XNOR2_X1 U1549 ( .A(n1354), .B(n1355), .ZN(p11_S[65]) );
  OAI221_X1 U1707 ( .B1(reg2[4]), .B2(n1403), .C1(n2817), .C2(n1404), .A(n1530), .ZN(n1511) );
  AOI22_X1 U1706 ( .A1(reg2[3]), .A2(n1323), .B1(n1324), .B2(
        p11_minus_A_shifted_16_), .ZN(n1529) );
  OAI221_X1 U1705 ( .B1(reg2[2]), .B2(n1319), .C1(n2820), .C2(n1321), .A(n1529), .ZN(n1512) );
  OAI221_X1 U1702 ( .B1(reg2[6]), .B2(n1420), .C1(n2835), .C2(n1421), .A(n1527), .ZN(n1513) );
  AOI222_X1 U1692 ( .A1(n1511), .A2(n1512), .B1(n1511), .B2(n1513), .C1(n1512), 
        .C2(n1513), .ZN(n1360) );
  XNOR2_X1 U1704 ( .A(n1511), .B(n1512), .ZN(n1526) );
  XNOR2_X1 U1701 ( .A(n1526), .B(n1513), .ZN(n1508) );
  XNOR2_X1 U1709 ( .A(n1503), .B(n1531), .ZN(n1509) );
  NAND2_X1 U1891 ( .A1(A1[1]), .A2(n1657), .ZN(n1567) );
  NAND2_X1 U1893 ( .A1(A1[0]), .A2(A1[1]), .ZN(n1590) );
  OAI21_X1 U1750 ( .B1(reg2[12]), .B2(n1567), .A(n1568), .ZN(n1566) );
  NAND2_X1 U1749 ( .A1(n1566), .A2(p11_muxs_out_1__13_), .ZN(n1523) );
  XNOR2_X1 U1727 ( .A(p11_muxs_out_3__14_), .B(p11_muxs_out_2__14_), .ZN(n1547) );
  OAI222_X1 U1699 ( .A1(n1523), .A2(n1524), .B1(n1523), .B2(n1525), .C1(n1524), 
        .C2(n1525), .ZN(n1510) );
  AOI222_X1 U1691 ( .A1(n1508), .A2(n1509), .B1(n1508), .B2(n1510), .C1(n1509), 
        .C2(n1510), .ZN(n1359) );
  XNOR2_X1 U1683 ( .A(n1491), .B(n1492), .ZN(n1496) );
  AOI222_X1 U1673 ( .A1(n1360), .A2(n1359), .B1(n1360), .B2(n1361), .C1(n1359), 
        .C2(n1361), .ZN(p11_C[64]) );
  XNOR2_X1 U1551 ( .A(n1358), .B(n1359), .ZN(p11_S[64]) );
  XNOR2_X1 U1700 ( .A(n1509), .B(n1508), .ZN(n1522) );
  XNOR2_X1 U1723 ( .A(n1524), .B(n1525), .ZN(n1546) );
  OAI221_X1 U1754 ( .B1(reg2[4]), .B2(n1420), .C1(n2817), .C2(n1421), .A(n1571), .ZN(n1554) );
  AOI222_X1 U1738 ( .A1(p11_muxs_out_2__13_), .A2(p11_muxs_out_3__13_), .B1(
        p11_muxs_out_2__13_), .B2(n1554), .C1(p11_muxs_out_3__13_), .C2(n1554), 
        .ZN(n1516) );
  AOI22_X1 U1735 ( .A1(reg2[1]), .A2(n1321), .B1(n1319), .B2(
        p11_minus_A_shifted_14_), .ZN(n1552) );
  AOI221_X1 U1734 ( .B1(n1323), .B2(reg2[2]), .C1(n1324), .C2(n2820), .A(n1552), .ZN(n1517) );
  XNOR2_X1 U1733 ( .A(n1516), .B(n1517), .ZN(n1550) );
  OAI221_X1 U1731 ( .B1(reg2[3]), .B2(n1403), .C1(p11_minus_A_shifted_16_), 
        .C2(n1404), .A(n1551), .ZN(n1518) );
  XNOR2_X1 U1730 ( .A(n1550), .B(n1518), .ZN(n1520) );
  XNOR2_X1 U1753 ( .A(p11_muxs_out_3__13_), .B(n1554), .ZN(n1570) );
  OAI21_X1 U1748 ( .B1(n1566), .B2(p11_muxs_out_1__13_), .A(n1523), .ZN(n1544)
         );
  OAI222_X1 U1784 ( .A1(reg2[12]), .A2(n1590), .B1(n2863), .B2(n1591), .C1(
        reg2[11]), .C2(n1567), .ZN(n1589) );
  NAND2_X1 U1783 ( .A1(n1589), .A2(p11_muxs_out_1__12_), .ZN(n1545) );
  AOI222_X1 U1720 ( .A1(n1543), .A2(n1544), .B1(n1543), .B2(n1545), .C1(n1544), 
        .C2(n1545), .ZN(n1521) );
  AOI222_X1 U1697 ( .A1(n1519), .A2(n1520), .B1(n1519), .B2(n1521), .C1(n1520), 
        .C2(n1521), .ZN(n1365) );
  OAI222_X1 U1695 ( .A1(n1515), .A2(n1516), .B1(n1515), .B2(n1517), .C1(n1516), 
        .C2(n1517), .ZN(n1514) );
  AOI222_X1 U1693 ( .A1(n1364), .A2(n1365), .B1(n1364), .B2(n1362), .C1(n1365), 
        .C2(n1362), .ZN(p11_C[63]) );
  XNOR2_X1 U1553 ( .A(n1362), .B(n1363), .ZN(p11_S[63]) );
  XNOR2_X1 U1719 ( .A(n1542), .B(n1521), .ZN(n1368) );
  XNOR2_X1 U1746 ( .A(n1543), .B(n1565), .ZN(n1539) );
  OAI22_X1 U1761 ( .A1(n2838), .A2(n1326), .B1(n1409), .B2(reg2[0]), .ZN(n1574) );
  OAI221_X1 U1760 ( .B1(n1411), .B2(p11_minus_A_shifted_14_), .C1(n1412), .C2(
        reg2[1]), .A(n1574), .ZN(n1537) );
  OAI221_X1 U1758 ( .B1(reg2[2]), .B2(n1403), .C1(n2820), .C2(n1404), .A(n1573), .ZN(n1535) );
  XNOR2_X1 U1756 ( .A(n1538), .B(n1572), .ZN(n1540) );
  XNOR2_X1 U1776 ( .A(p11_muxs_out_2__12_), .B(n1586), .ZN(n1562) );
  OAI21_X1 U1782 ( .B1(n1589), .B2(p11_muxs_out_1__12_), .A(n1545), .ZN(n1563)
         );
  OAI21_X1 U1801 ( .B1(reg2[11]), .B2(n1590), .A(n1607), .ZN(n1588) );
  NAND2_X1 U1781 ( .A1(p11_muxs_out_1__11_), .A2(n1588), .ZN(n1564) );
  AOI222_X1 U1744 ( .A1(n1562), .A2(n1563), .B1(n1562), .B2(n1564), .C1(n1563), 
        .C2(n1564), .ZN(n1541) );
  AOI222_X1 U1718 ( .A1(n1539), .A2(n1540), .B1(n1539), .B2(n1541), .C1(n1540), 
        .C2(n1541), .ZN(n1369) );
  AOI222_X1 U1716 ( .A1(n1535), .A2(n1536), .B1(n1535), .B2(n1537), .C1(n1536), 
        .C2(n1537), .ZN(n1366) );
  AOI222_X1 U1715 ( .A1(n1368), .A2(n1369), .B1(n1368), .B2(n1366), .C1(n1369), 
        .C2(n1366), .ZN(p11_C[62]) );
  XNOR2_X1 U1555 ( .A(n1366), .B(n1367), .ZN(p11_S[62]) );
  XNOR2_X1 U1743 ( .A(n1561), .B(n1541), .ZN(n1372) );
  OAI221_X1 U1789 ( .B1(reg2[1]), .B2(n1403), .C1(p11_minus_A_shifted_14_), 
        .C2(n1404), .A(n1593), .ZN(n1555) );
  NOR2_X1 U1786 ( .A1(n1575), .A2(n2838), .ZN(n1592) );
  XNOR2_X1 U1780 ( .A(n1563), .B(n1564), .ZN(n1585) );
  XNOR2_X1 U1800 ( .A(n1588), .B(p11_muxs_out_1__11_), .ZN(n1594) );
  OAI21_X1 U1824 ( .B1(reg2[10]), .B2(n1590), .A(n1621), .ZN(n1620) );
  NAND2_X1 U1823 ( .A1(p11_muxs_out_1__10_), .A2(n1620), .ZN(n1596) );
  AOI222_X1 U1791 ( .A1(n1594), .A2(n1595), .B1(n1594), .B2(n1596), .C1(n1595), 
        .C2(n1596), .ZN(n1560) );
  AOI222_X1 U1742 ( .A1(n1558), .A2(n1559), .B1(n1558), .B2(n1560), .C1(n1559), 
        .C2(n1560), .ZN(n1373) );
  OAI221_X1 U1741 ( .B1(reg2[0]), .B2(n1412), .C1(n2838), .C2(n1411), .A(n1319), .ZN(n1556) );
  AOI222_X1 U1740 ( .A1(n1555), .A2(A1[13]), .B1(n1555), .B2(n1556), .C1(
        A1[13]), .C2(n1556), .ZN(n1370) );
  AOI222_X1 U1739 ( .A1(n1372), .A2(n1373), .B1(n1372), .B2(n1370), .C1(n1373), 
        .C2(n1370), .ZN(p11_C[61]) );
  XNOR2_X1 U1557 ( .A(n1370), .B(n1371), .ZN(p11_S[61]) );
  OAI221_X1 U1810 ( .B1(reg2[0]), .B2(n1403), .C1(n2838), .C2(n1404), .A(n1612), .ZN(n1597) );
  OAI221_X1 U1807 ( .B1(reg2[2]), .B2(n1420), .C1(n2820), .C2(n1421), .A(n1611), .ZN(n1598) );
  XNOR2_X1 U1806 ( .A(n1610), .B(n1598), .ZN(n1581) );
  AOI22_X1 U1803 ( .A1(p11_muxs_out_2__11_), .A2(n1609), .B1(n1596), .B2(n1595), .ZN(n1606) );
  XNOR2_X1 U1799 ( .A(n1606), .B(n1594), .ZN(n1582) );
  OAI21_X1 U1822 ( .B1(p11_muxs_out_1__10_), .B2(n1620), .A(n1596), .ZN(n1616)
         );
  AOI222_X1 U1816 ( .A1(n1614), .A2(n1615), .B1(n1614), .B2(n1616), .C1(n1615), 
        .C2(n1616), .ZN(n1583) );
  AOI222_X1 U1772 ( .A1(n1581), .A2(n1582), .B1(n1581), .B2(n1583), .C1(n1582), 
        .C2(n1583), .ZN(n1374) );
  OAI221_X1 U1833 ( .B1(reg2[1]), .B2(n1420), .C1(p11_minus_A_shifted_14_), 
        .C2(n1421), .A(n1622), .ZN(n1600) );
  NOR2_X1 U1830 ( .A1(n1613), .A2(n2838), .ZN(n1601) );
  XNOR2_X1 U1797 ( .A(n1583), .B(n1605), .ZN(n1380) );
  NOR2_X1 U1848 ( .A1(reg2[8]), .A2(n1567), .ZN(n1637) );
  AOI222_X1 U1835 ( .A1(n1623), .A2(n1624), .B1(n1623), .B2(n1625), .C1(n1624), 
        .C2(n1625), .ZN(n1604) );
  AOI22_X1 U1849 ( .A1(p11_muxs_out_1__9_), .A2(p11_muxs_out_2__9_), .B1(n1624), .B2(n1623), .ZN(n1636) );
  XNOR2_X1 U1846 ( .A(n1636), .B(n1625), .ZN(n1626) );
  AOI22_X1 U1845 ( .A1(reg2[0]), .A2(n1421), .B1(n1420), .B2(n2838), .ZN(n1635) );
  OAI221_X1 U1843 ( .B1(n1632), .B2(p11_minus_A_shifted_14_), .C1(n1633), .C2(
        reg2[1]), .A(n1634), .ZN(n1617) );
  OAI21_X1 U1869 ( .B1(reg2[7]), .B2(n1567), .A(n1647), .ZN(n1631) );
  AOI222_X1 U1840 ( .A1(p11_muxs_out_1__8_), .A2(p11_muxs_out_2__8_), .B1(
        p11_muxs_out_1__8_), .B2(n1631), .C1(p11_muxs_out_2__8_), .C2(n1631), 
        .ZN(n1629) );
  NAND2_X1 U1818 ( .A1(p11_muxs_out_3__9_), .A2(n1617), .ZN(n1382) );
  XNOR2_X1 U1841 ( .A(n1626), .B(n1627), .ZN(n1630) );
  XNOR2_X1 U1839 ( .A(n1630), .B(n1629), .ZN(n1386) );
  AOI22_X1 U1882 ( .A1(reg2[7]), .A2(n1591), .B1(n1590), .B2(n2831), .ZN(n1653) );
  NOR2_X1 U1890 ( .A1(reg2[5]), .A2(n1567), .ZN(n1656) );
  NOR2_X1 U1876 ( .A1(n1649), .A2(n1650), .ZN(n1642) );
  XNOR2_X1 U1888 ( .A(p11_muxs_out_1__6_), .B(n1649), .ZN(n1655) );
  NAND2_X1 U1887 ( .A1(n1655), .A2(p11_muxs_out_2__6_), .ZN(n1398) );
  AOI222_X1 U1872 ( .A1(n1396), .A2(n1399), .B1(n1396), .B2(n1398), .C1(n1399), 
        .C2(n1398), .ZN(p11_C[55]) );
  AOI22_X1 U1571 ( .A1(p11_muxs_out_3__7_), .A2(n1397), .B1(n1398), .B2(n1399), 
        .ZN(n1395) );
  XNOR2_X1 U1570 ( .A(n1395), .B(n1396), .ZN(p11_S[55]) );
  OAI21_X1 U1886 ( .B1(n1655), .B2(p11_muxs_out_2__6_), .A(n1398), .ZN(n1400)
         );
  NOR2_X1 U1885 ( .A1(n1654), .A2(n1400), .ZN(p11_C[54]) );
  XNOR2_X1 U1573 ( .A(p11_muxs_out_3__6_), .B(n1400), .ZN(p11_S[54]) );
  AOI222_X1 U1838 ( .A1(n1388), .A2(n1389), .B1(n1388), .B2(n1386), .C1(n1389), 
        .C2(n1386), .ZN(p11_C[57]) );
  AOI222_X1 U1793 ( .A1(n1380), .A2(n1381), .B1(n1380), .B2(n1378), .C1(n1381), 
        .C2(n1378), .ZN(p11_C[59]) );
  AOI21_X1 U2133 ( .B1(n1918), .B2(n1919), .A(n1665), .ZN(n1916) );
  AOI22_X1 U2154 ( .A1(A2[11]), .A2(n1919), .B1(A2[12]), .B2(n1918), .ZN(n1915) );
  AOI22_X1 U1899 ( .A1(reg4[13]), .A2(n1662), .B1(n1663), .B2(n2859), .ZN(
        n1661) );
  OAI221_X1 U1898 ( .B1(reg4[12]), .B2(n1658), .C1(n2858), .C2(n1660), .A(
        n1661), .ZN(p10_final_product2_26_) );
  AOI22_X1 U1942 ( .A1(reg4[12]), .A2(n1662), .B1(n1663), .B2(n2858), .ZN(
        n1742) );
  AOI22_X1 U1957 ( .A1(reg4[12]), .A2(n1746), .B1(n1747), .B2(n2858), .ZN(
        n1763) );
  OAI221_X1 U1956 ( .B1(reg4[11]), .B2(n1743), .C1(n2861), .C2(n1744), .A(
        n1763), .ZN(n1753) );
  OAI221_X1 U1955 ( .B1(reg4[13]), .B2(n1760), .C1(n2859), .C2(n1761), .A(
        n1762), .ZN(n1756) );
  AOI22_X1 U1953 ( .A1(reg4[10]), .A2(n1662), .B1(n1663), .B2(n2810), .ZN(
        n1759) );
  OAI221_X1 U1952 ( .B1(reg4[9]), .B2(n1658), .C1(n2814), .C2(n1660), .A(n1759), .ZN(n1755) );
  AOI222_X1 U1948 ( .A1(n1753), .A2(n1754), .B1(n1753), .B2(n1755), .C1(n1754), 
        .C2(n1755), .ZN(n1669) );
  AOI22_X1 U1947 ( .A1(reg4[11]), .A2(n1751), .B1(n1752), .B2(n2861), .ZN(
        n1750) );
  AOI221_X1 U1946 ( .B1(reg4[10]), .B2(n1665), .C1(n2810), .C2(n1749), .A(
        n1750), .ZN(n1670) );
  AOI22_X1 U1945 ( .A1(reg4[13]), .A2(n1746), .B1(n1747), .B2(n2859), .ZN(
        n1745) );
  OAI221_X1 U1944 ( .B1(reg4[12]), .B2(n1743), .C1(n2858), .C2(n1744), .A(
        n1745), .ZN(n1667) );
  AOI222_X1 U1943 ( .A1(n1669), .A2(n1670), .B1(n1669), .B2(n1667), .C1(n1670), 
        .C2(n1667), .ZN(p10_C[71]) );
  XNOR2_X1 U1903 ( .A(n1667), .B(n1668), .ZN(p10_S[71]) );
  OAI221_X1 U1966 ( .B1(reg4[12]), .B2(n1760), .C1(n2858), .C2(n1761), .A(
        n1762), .ZN(n1673) );
  AOI22_X1 U1965 ( .A1(reg4[11]), .A2(n1746), .B1(n1747), .B2(n2861), .ZN(
        n1768) );
  OAI221_X1 U1964 ( .B1(reg4[10]), .B2(n1743), .C1(n2810), .C2(n1744), .A(
        n1768), .ZN(n1764) );
  OAI221_X1 U1987 ( .B1(reg4[11]), .B2(n1760), .C1(n2861), .C2(n1761), .A(
        n1790), .ZN(n1771) );
  AOI22_X1 U1985 ( .A1(reg4[10]), .A2(n1746), .B1(n1747), .B2(n2810), .ZN(
        n1789) );
  OAI221_X1 U1984 ( .B1(reg4[9]), .B2(n1743), .C1(n2814), .C2(n1744), .A(n1789), .ZN(n1772) );
  AOI222_X1 U1968 ( .A1(n1771), .A2(n1772), .B1(n1771), .B2(n1773), .C1(n1772), 
        .C2(n1773), .ZN(n1766) );
  AOI222_X1 U1958 ( .A1(n1764), .A2(n1676), .B1(n1764), .B2(n1765), .C1(n1676), 
        .C2(n1765), .ZN(n1672) );
  XNOR2_X1 U1954 ( .A(n1753), .B(n1756), .ZN(n1757) );
  XNOR2_X1 U1951 ( .A(n1757), .B(n1755), .ZN(n1675) );
  AOI222_X1 U1950 ( .A1(n1676), .A2(n1672), .B1(n1676), .B2(n1675), .C1(n1672), 
        .C2(n1675), .ZN(p10_C[70]) );
  AOI22_X1 U1906 ( .A1(n1673), .A2(n1674), .B1(n1675), .B2(n1676), .ZN(n1671)
         );
  XNOR2_X1 U1905 ( .A(n1671), .B(n1672), .ZN(p10_S[70]) );
  XNOR2_X1 U1986 ( .A(p10_muxs_out_3__20_), .B(n1771), .ZN(n1788) );
  AOI22_X1 U1982 ( .A1(reg4[8]), .A2(n1662), .B1(n1663), .B2(n2832), .ZN(n1787) );
  OAI221_X1 U1981 ( .B1(reg4[7]), .B2(n1658), .C1(n2830), .C2(n1660), .A(n1787), .ZN(n1777) );
  AOI22_X1 U1996 ( .A1(reg4[8]), .A2(n1744), .B1(n1743), .B2(n2832), .ZN(n1798) );
  AOI221_X1 U1995 ( .B1(n1746), .B2(reg4[9]), .C1(n1747), .C2(n2814), .A(n1798), .ZN(n1783) );
  OAI221_X1 U1998 ( .B1(reg4[10]), .B2(n1760), .C1(n2810), .C2(n1761), .A(
        n1799), .ZN(n1785) );
  AOI222_X1 U1978 ( .A1(p10_muxs_out_3__19_), .A2(n1783), .B1(
        p10_muxs_out_3__19_), .B2(n1784), .C1(n1783), .C2(n1784), .ZN(n1778)
         );
  AOI222_X1 U1972 ( .A1(n1776), .A2(n1777), .B1(n1776), .B2(n1778), .C1(n1777), 
        .C2(n1778), .ZN(n1679) );
  AOI22_X1 U1971 ( .A1(reg4[9]), .A2(n1751), .B1(n1752), .B2(n2814), .ZN(n1775) );
  AOI221_X1 U1970 ( .B1(reg4[8]), .B2(n1665), .C1(n2832), .C2(n1749), .A(n1775), .ZN(n1680) );
  XNOR2_X1 U1962 ( .A(n1766), .B(n1767), .ZN(n1677) );
  AOI222_X1 U1961 ( .A1(n1679), .A2(n1680), .B1(n1679), .B2(n1677), .C1(n1680), 
        .C2(n1677), .ZN(p10_C[69]) );
  XNOR2_X1 U1908 ( .A(n1677), .B(n1678), .ZN(p10_S[69]) );
  XNOR2_X1 U1977 ( .A(n1782), .B(n1778), .ZN(n1681) );
  XNOR2_X1 U1997 ( .A(p10_muxs_out_3__19_), .B(n1785), .ZN(n1797) );
  AOI22_X1 U2015 ( .A1(reg4[8]), .A2(n1746), .B1(n1747), .B2(n2832), .ZN(n1813) );
  OAI221_X1 U2014 ( .B1(reg4[7]), .B2(n1743), .C1(n2830), .C2(n1744), .A(n1813), .ZN(n1802) );
  AOI22_X1 U2012 ( .A1(reg4[6]), .A2(n1662), .B1(n1663), .B2(n2815), .ZN(n1812) );
  OAI221_X1 U2011 ( .B1(reg4[5]), .B2(n1658), .C1(n2813), .C2(n1660), .A(n1812), .ZN(n1803) );
  AOI222_X1 U2003 ( .A1(p10_muxs_out_2__17_), .A2(n1802), .B1(
        p10_muxs_out_2__17_), .B2(n1803), .C1(n1802), .C2(n1803), .ZN(n1780)
         );
  OAI221_X1 U2018 ( .B1(reg4[9]), .B2(n1760), .C1(n2814), .C2(n1761), .A(n1815), .ZN(n1800) );
  AOI222_X1 U2001 ( .A1(p10_muxs_out_3__18_), .A2(n1800), .B1(
        p10_muxs_out_3__18_), .B2(n1801), .C1(n1800), .C2(n1801), .ZN(n1781)
         );
  OAI222_X1 U1975 ( .A1(n1779), .A2(n1780), .B1(n1779), .B2(n1781), .C1(n1780), 
        .C2(n1781), .ZN(n1683) );
  AOI222_X1 U1973 ( .A1(n1681), .A2(n1685), .B1(n1681), .B2(n1684), .C1(n1685), 
        .C2(n1684), .ZN(p10_C[68]) );
  AOI22_X1 U1911 ( .A1(p10_muxs_out_3__19_), .A2(n1683), .B1(n1684), .B2(n1685), .ZN(n1682) );
  XNOR2_X1 U1910 ( .A(n1681), .B(n1682), .ZN(p10_S[68]) );
  XNOR2_X1 U2000 ( .A(n1780), .B(n1781), .ZN(n1796) );
  XNOR2_X1 U1993 ( .A(n1796), .B(n1779), .ZN(n1686) );
  XNOR2_X1 U2013 ( .A(p10_muxs_out_2__17_), .B(n1802), .ZN(n1810) );
  XNOR2_X1 U2010 ( .A(n1810), .B(n1803), .ZN(n1793) );
  AOI222_X1 U2036 ( .A1(p10_muxs_out_2__16_), .A2(p10_muxs_out_3__16_), .B1(
        p10_muxs_out_2__16_), .B2(n1830), .C1(p10_muxs_out_3__16_), .C2(n1830), 
        .ZN(n1809) );
  AOI222_X1 U2008 ( .A1(p10_muxs_out_2__17_), .A2(n1808), .B1(
        p10_muxs_out_2__17_), .B2(n1809), .C1(n1808), .C2(n1809), .ZN(n1794)
         );
  XNOR2_X1 U2016 ( .A(p10_muxs_out_2__18_), .B(n1814), .ZN(n1795) );
  AOI222_X1 U1992 ( .A1(n1793), .A2(n1794), .B1(n1793), .B2(n1795), .C1(n1794), 
        .C2(n1795), .ZN(n1689) );
  OAI22_X1 U1991 ( .A1(n2830), .A2(n1751), .B1(n1752), .B2(reg4[7]), .ZN(n1792) );
  AOI221_X1 U1990 ( .B1(n2815), .B2(n1749), .C1(reg4[6]), .C2(n1665), .A(n1792), .ZN(n1688) );
  AOI222_X1 U1989 ( .A1(n1686), .A2(n1689), .B1(n1686), .B2(n1688), .C1(n1689), 
        .C2(n1688), .ZN(p10_C[67]) );
  XNOR2_X1 U1913 ( .A(n1688), .B(n1689), .ZN(n1687) );
  AOI22_X1 U2033 ( .A1(reg4[7]), .A2(n1746), .B1(n1747), .B2(n2830), .ZN(n1828) );
  OAI221_X1 U2032 ( .B1(reg4[6]), .B2(n1743), .C1(n2815), .C2(n1744), .A(n1828), .ZN(n1804) );
  AOI22_X1 U2031 ( .A1(reg4[5]), .A2(n1662), .B1(n1663), .B2(n2813), .ZN(n1827) );
  OAI221_X1 U2030 ( .B1(reg4[4]), .B2(n1658), .C1(n2818), .C2(n1660), .A(n1827), .ZN(n1805) );
  XNOR2_X1 U2029 ( .A(n1804), .B(n1805), .ZN(n1824) );
  OAI221_X1 U2027 ( .B1(reg4[8]), .B2(n1760), .C1(n2832), .C2(n1761), .A(n1825), .ZN(n1806) );
  XNOR2_X1 U2026 ( .A(n1824), .B(n1806), .ZN(n1816) );
  XNOR2_X1 U2047 ( .A(p10_muxs_out_3__16_), .B(p10_muxs_out_2__16_), .ZN(n1839) );
  XNOR2_X1 U2046 ( .A(n1839), .B(p10_muxs_out_1__16_), .ZN(n1820) );
  AOI222_X1 U2043 ( .A1(p10_muxs_out_3__15_), .A2(p10_muxs_out_2__15_), .B1(
        p10_muxs_out_3__15_), .B2(n1838), .C1(p10_muxs_out_2__15_), .C2(n1838), 
        .ZN(n1821) );
  OAI221_X1 U2048 ( .B1(reg4[7]), .B2(n1760), .C1(n2830), .C2(n1761), .A(n1840), .ZN(n1823) );
  AOI222_X1 U2023 ( .A1(n1820), .A2(n1821), .B1(n1820), .B2(n1822), .C1(n1821), 
        .C2(n1822), .ZN(n1818) );
  AOI222_X1 U2020 ( .A1(n1816), .A2(n1817), .B1(n1816), .B2(n1818), .C1(n1817), 
        .C2(n1818), .ZN(n1692) );
  XNOR2_X1 U2006 ( .A(n1795), .B(n1807), .ZN(n1693) );
  AOI222_X1 U2005 ( .A1(n1804), .A2(n1805), .B1(n1804), .B2(n1806), .C1(n1805), 
        .C2(n1806), .ZN(n1690) );
  AOI222_X1 U2004 ( .A1(n1692), .A2(n1693), .B1(n1692), .B2(n1690), .C1(n1693), 
        .C2(n1690), .ZN(p10_C[66]) );
  XNOR2_X1 U1914 ( .A(n1690), .B(n1691), .ZN(p10_S[66]) );
  AOI22_X1 U2057 ( .A1(reg4[6]), .A2(n1746), .B1(n1747), .B2(n2815), .ZN(n1847) );
  OAI221_X1 U2056 ( .B1(reg4[5]), .B2(n1743), .C1(n2813), .C2(n1744), .A(n1847), .ZN(n1834) );
  AOI22_X1 U2054 ( .A1(reg4[4]), .A2(n1662), .B1(n1663), .B2(n2818), .ZN(n1846) );
  OAI221_X1 U2053 ( .B1(reg4[3]), .B2(n1658), .C1(p10_minus_A_shifted_16_), 
        .C2(n1660), .A(n1846), .ZN(n1835) );
  AOI222_X1 U2039 ( .A1(p10_muxs_out_1__15_), .A2(n1834), .B1(
        p10_muxs_out_1__15_), .B2(n1835), .C1(n1834), .C2(n1835), .ZN(n1696)
         );
  XNOR2_X1 U2055 ( .A(p10_muxs_out_1__15_), .B(n1834), .ZN(n1844) );
  XNOR2_X1 U2052 ( .A(n1844), .B(n1835), .ZN(n1831) );
  NOR2_X1 U2080 ( .A1(p10_muxs_out_1__14_), .A2(n1873), .ZN(n1841) );
  XNOR2_X1 U2079 ( .A(p10_muxs_out_1__15_), .B(p10_muxs_out_3__15_), .ZN(n1872) );
  XNOR2_X1 U2078 ( .A(n1872), .B(p10_muxs_out_2__15_), .ZN(n1842) );
  OAI221_X1 U2092 ( .B1(reg4[5]), .B2(n1760), .C1(n2813), .C2(n1761), .A(n1888), .ZN(n1874) );
  AOI222_X1 U2081 ( .A1(p10_muxs_out_3__14_), .A2(p10_muxs_out_2__14_), .B1(
        p10_muxs_out_3__14_), .B2(n1874), .C1(p10_muxs_out_2__14_), .C2(n1874), 
        .ZN(n1843) );
  AOI222_X1 U2051 ( .A1(n1841), .A2(n1842), .B1(n1841), .B2(n1843), .C1(n1842), 
        .C2(n1843), .ZN(n1832) );
  XNOR2_X1 U2045 ( .A(n1823), .B(n1820), .ZN(n1837) );
  XNOR2_X1 U2042 ( .A(n1837), .B(n1821), .ZN(n1833) );
  AOI222_X1 U2038 ( .A1(n1831), .A2(n1832), .B1(n1831), .B2(n1833), .C1(n1832), 
        .C2(n1833), .ZN(n1697) );
  XNOR2_X1 U2022 ( .A(n1819), .B(n1818), .ZN(n1694) );
  AOI222_X1 U2021 ( .A1(n1696), .A2(n1697), .B1(n1696), .B2(n1694), .C1(n1697), 
        .C2(n1694), .ZN(p10_C[65]) );
  XNOR2_X1 U1916 ( .A(n1694), .B(n1695), .ZN(p10_S[65]) );
  AOI22_X1 U2075 ( .A1(reg4[5]), .A2(n1746), .B1(n1747), .B2(n2813), .ZN(n1870) );
  OAI221_X1 U2074 ( .B1(reg4[4]), .B2(n1743), .C1(n2818), .C2(n1744), .A(n1870), .ZN(n1851) );
  AOI22_X1 U2073 ( .A1(reg4[3]), .A2(n1662), .B1(n1663), .B2(
        p10_minus_A_shifted_16_), .ZN(n1869) );
  OAI221_X1 U2072 ( .B1(reg4[2]), .B2(n1658), .C1(n2821), .C2(n1660), .A(n1869), .ZN(n1852) );
  OAI221_X1 U2069 ( .B1(reg4[6]), .B2(n1760), .C1(n2815), .C2(n1761), .A(n1867), .ZN(n1853) );
  AOI222_X1 U2059 ( .A1(n1851), .A2(n1852), .B1(n1851), .B2(n1853), .C1(n1852), 
        .C2(n1853), .ZN(n1700) );
  XNOR2_X1 U2071 ( .A(n1851), .B(n1852), .ZN(n1866) );
  XNOR2_X1 U2068 ( .A(n1866), .B(n1853), .ZN(n1848) );
  XNOR2_X1 U2076 ( .A(n1843), .B(n1871), .ZN(n1849) );
  NAND2_X1 U2258 ( .A1(A2[1]), .A2(n1997), .ZN(n1907) );
  NAND2_X1 U2260 ( .A1(A2[0]), .A2(A2[1]), .ZN(n1930) );
  OAI21_X1 U2117 ( .B1(reg4[12]), .B2(n1907), .A(n1908), .ZN(n1906) );
  NAND2_X1 U2116 ( .A1(n1906), .A2(p10_muxs_out_1__13_), .ZN(n1863) );
  XNOR2_X1 U2094 ( .A(p10_muxs_out_3__14_), .B(p10_muxs_out_2__14_), .ZN(n1887) );
  OAI222_X1 U2066 ( .A1(n1863), .A2(n1864), .B1(n1863), .B2(n1865), .C1(n1864), 
        .C2(n1865), .ZN(n1850) );
  AOI222_X1 U2058 ( .A1(n1848), .A2(n1849), .B1(n1848), .B2(n1850), .C1(n1849), 
        .C2(n1850), .ZN(n1699) );
  XNOR2_X1 U2050 ( .A(n1831), .B(n1832), .ZN(n1836) );
  AOI222_X1 U2040 ( .A1(n1700), .A2(n1699), .B1(n1700), .B2(n1701), .C1(n1699), 
        .C2(n1701), .ZN(p10_C[64]) );
  XNOR2_X1 U1918 ( .A(n1698), .B(n1699), .ZN(p10_S[64]) );
  XNOR2_X1 U2067 ( .A(n1849), .B(n1848), .ZN(n1862) );
  XNOR2_X1 U2090 ( .A(n1864), .B(n1865), .ZN(n1886) );
  OAI221_X1 U2121 ( .B1(reg4[4]), .B2(n1760), .C1(n2818), .C2(n1761), .A(n1911), .ZN(n1894) );
  AOI222_X1 U2105 ( .A1(p10_muxs_out_2__13_), .A2(p10_muxs_out_3__13_), .B1(
        p10_muxs_out_2__13_), .B2(n1894), .C1(p10_muxs_out_3__13_), .C2(n1894), 
        .ZN(n1856) );
  AOI22_X1 U2102 ( .A1(reg4[1]), .A2(n1660), .B1(n1658), .B2(
        p10_minus_A_shifted_14_), .ZN(n1892) );
  AOI221_X1 U2101 ( .B1(n1662), .B2(reg4[2]), .C1(n1663), .C2(n2821), .A(n1892), .ZN(n1857) );
  XNOR2_X1 U2100 ( .A(n1856), .B(n1857), .ZN(n1890) );
  AOI22_X1 U2099 ( .A1(reg4[4]), .A2(n1746), .B1(n1747), .B2(n2818), .ZN(n1891) );
  OAI221_X1 U2098 ( .B1(reg4[3]), .B2(n1743), .C1(p10_minus_A_shifted_16_), 
        .C2(n1744), .A(n1891), .ZN(n1858) );
  XNOR2_X1 U2097 ( .A(n1890), .B(n1858), .ZN(n1860) );
  XNOR2_X1 U2120 ( .A(p10_muxs_out_3__13_), .B(n1894), .ZN(n1910) );
  OAI21_X1 U2115 ( .B1(n1906), .B2(p10_muxs_out_1__13_), .A(n1863), .ZN(n1884)
         );
  OAI222_X1 U2151 ( .A1(reg4[12]), .A2(n1930), .B1(n2858), .B2(n1931), .C1(
        reg4[11]), .C2(n1907), .ZN(n1929) );
  NAND2_X1 U2150 ( .A1(n1929), .A2(p10_muxs_out_1__12_), .ZN(n1885) );
  AOI222_X1 U2087 ( .A1(n1883), .A2(n1884), .B1(n1883), .B2(n1885), .C1(n1884), 
        .C2(n1885), .ZN(n1861) );
  AOI222_X1 U2064 ( .A1(n1859), .A2(n1860), .B1(n1859), .B2(n1861), .C1(n1860), 
        .C2(n1861), .ZN(n1705) );
  OAI222_X1 U2062 ( .A1(n1855), .A2(n1856), .B1(n1855), .B2(n1857), .C1(n1856), 
        .C2(n1857), .ZN(n1854) );
  AOI222_X1 U2060 ( .A1(n1704), .A2(n1705), .B1(n1704), .B2(n1702), .C1(n1705), 
        .C2(n1702), .ZN(p10_C[63]) );
  XNOR2_X1 U1920 ( .A(n1702), .B(n1703), .ZN(p10_S[63]) );
  XNOR2_X1 U2086 ( .A(n1882), .B(n1861), .ZN(n1708) );
  XNOR2_X1 U2113 ( .A(n1883), .B(n1905), .ZN(n1879) );
  OAI22_X1 U2128 ( .A1(n2839), .A2(n1665), .B1(n1749), .B2(reg4[0]), .ZN(n1914) );
  OAI221_X1 U2127 ( .B1(n1751), .B2(p10_minus_A_shifted_14_), .C1(n1752), .C2(
        reg4[1]), .A(n1914), .ZN(n1877) );
  AOI22_X1 U2126 ( .A1(reg4[3]), .A2(n1746), .B1(n1747), .B2(
        p10_minus_A_shifted_16_), .ZN(n1913) );
  OAI221_X1 U2125 ( .B1(reg4[2]), .B2(n1743), .C1(n2821), .C2(n1744), .A(n1913), .ZN(n1875) );
  XNOR2_X1 U2123 ( .A(n1878), .B(n1912), .ZN(n1880) );
  OAI21_X1 U2149 ( .B1(n1929), .B2(p10_muxs_out_1__12_), .A(n1885), .ZN(n1903)
         );
  OAI21_X1 U2168 ( .B1(reg4[11]), .B2(n1930), .A(n1947), .ZN(n1928) );
  NAND2_X1 U2148 ( .A1(p10_muxs_out_1__11_), .A2(n1928), .ZN(n1904) );
  AOI222_X1 U2111 ( .A1(n1902), .A2(n1903), .B1(n1902), .B2(n1904), .C1(n1903), 
        .C2(n1904), .ZN(n1881) );
  AOI222_X1 U2085 ( .A1(n1879), .A2(n1880), .B1(n1879), .B2(n1881), .C1(n1880), 
        .C2(n1881), .ZN(n1709) );
  AOI222_X1 U2083 ( .A1(n1875), .A2(n1876), .B1(n1875), .B2(n1877), .C1(n1876), 
        .C2(n1877), .ZN(n1706) );
  AOI222_X1 U2082 ( .A1(n1708), .A2(n1709), .B1(n1708), .B2(n1706), .C1(n1709), 
        .C2(n1706), .ZN(p10_C[62]) );
  XNOR2_X1 U1922 ( .A(n1706), .B(n1707), .ZN(p10_S[62]) );
  XNOR2_X1 U2110 ( .A(n1901), .B(n1881), .ZN(n1712) );
  AOI22_X1 U2157 ( .A1(reg4[2]), .A2(n1746), .B1(n1747), .B2(n2821), .ZN(n1933) );
  OAI221_X1 U2156 ( .B1(reg4[1]), .B2(n1743), .C1(p10_minus_A_shifted_14_), 
        .C2(n1744), .A(n1933), .ZN(n1895) );
  NOR2_X1 U2153 ( .A1(n1915), .A2(n2839), .ZN(n1932) );
  XNOR2_X1 U2167 ( .A(n1928), .B(p10_muxs_out_1__11_), .ZN(n1934) );
  OAI21_X1 U2191 ( .B1(reg4[10]), .B2(n1930), .A(n1961), .ZN(n1960) );
  NAND2_X1 U2190 ( .A1(p10_muxs_out_1__10_), .A2(n1960), .ZN(n1936) );
  AOI222_X1 U2158 ( .A1(n1934), .A2(n1935), .B1(n1934), .B2(n1936), .C1(n1935), 
        .C2(n1936), .ZN(n1900) );
  OAI221_X1 U2108 ( .B1(reg4[0]), .B2(n1752), .C1(n2839), .C2(n1751), .A(n1658), .ZN(n1896) );
  AOI222_X1 U2107 ( .A1(n1895), .A2(A2[13]), .B1(n1895), .B2(n1896), .C1(
        A2[13]), .C2(n1896), .ZN(n1710) );
  AOI222_X1 U2106 ( .A1(n1712), .A2(n1713), .B1(n1712), .B2(n1710), .C1(n1713), 
        .C2(n1710), .ZN(p10_C[61]) );
  XNOR2_X1 U1924 ( .A(n1710), .B(n1711), .ZN(p10_S[61]) );
  AOI22_X1 U2178 ( .A1(reg4[1]), .A2(n1746), .B1(n1747), .B2(
        p10_minus_A_shifted_14_), .ZN(n1952) );
  OAI221_X1 U2177 ( .B1(reg4[0]), .B2(n1743), .C1(n2839), .C2(n1744), .A(n1952), .ZN(n1937) );
  OAI221_X1 U2174 ( .B1(reg4[2]), .B2(n1760), .C1(n2821), .C2(n1761), .A(n1951), .ZN(n1938) );
  AOI222_X1 U2159 ( .A1(n1937), .A2(p10_muxs_out_3__11_), .B1(n1937), .B2(
        n1938), .C1(p10_muxs_out_3__11_), .C2(n1938), .ZN(n1716) );
  XNOR2_X1 U2176 ( .A(n1937), .B(p10_muxs_out_3__11_), .ZN(n1950) );
  XNOR2_X1 U2173 ( .A(n1950), .B(n1938), .ZN(n1921) );
  AOI22_X1 U2170 ( .A1(p10_muxs_out_2__11_), .A2(n1949), .B1(n1936), .B2(n1935), .ZN(n1946) );
  XNOR2_X1 U2166 ( .A(n1946), .B(n1934), .ZN(n1922) );
  OAI21_X1 U2189 ( .B1(p10_muxs_out_1__10_), .B2(n1960), .A(n1936), .ZN(n1956)
         );
  AOI222_X1 U2183 ( .A1(n1954), .A2(n1955), .B1(n1954), .B2(n1956), .C1(n1955), 
        .C2(n1956), .ZN(n1923) );
  AOI222_X1 U2139 ( .A1(n1921), .A2(n1922), .B1(n1921), .B2(n1923), .C1(n1922), 
        .C2(n1923), .ZN(n1714) );
  OAI221_X1 U2200 ( .B1(reg4[1]), .B2(n1760), .C1(p10_minus_A_shifted_14_), 
        .C2(n1761), .A(n1962), .ZN(n1940) );
  NOR2_X1 U2197 ( .A1(n1953), .A2(n2839), .ZN(n1941) );
  NOR2_X1 U2215 ( .A1(reg4[8]), .A2(n1907), .ZN(n1977) );
  AOI222_X1 U2202 ( .A1(n1963), .A2(n1964), .B1(n1963), .B2(n1965), .C1(n1964), 
        .C2(n1965), .ZN(n1944) );
  AOI22_X1 U2216 ( .A1(p10_muxs_out_1__9_), .A2(p10_muxs_out_2__9_), .B1(n1964), .B2(n1963), .ZN(n1976) );
  XNOR2_X1 U2213 ( .A(n1976), .B(n1965), .ZN(n1966) );
  AOI22_X1 U2212 ( .A1(reg4[0]), .A2(n1761), .B1(n1760), .B2(n2839), .ZN(n1975) );
  OAI221_X1 U2210 ( .B1(n1972), .B2(p10_minus_A_shifted_14_), .C1(n1973), .C2(
        reg4[1]), .A(n1974), .ZN(n1957) );
  OAI21_X1 U2236 ( .B1(reg4[7]), .B2(n1907), .A(n1987), .ZN(n1971) );
  AOI222_X1 U2203 ( .A1(n1966), .A2(n1967), .B1(n1966), .B2(n1968), .C1(n1967), 
        .C2(n1968), .ZN(n1724) );
  NAND2_X1 U2185 ( .A1(p10_muxs_out_3__9_), .A2(n1957), .ZN(n1722) );
  XNOR2_X1 U2208 ( .A(n1966), .B(n1967), .ZN(n1970) );
  XNOR2_X1 U2206 ( .A(n1970), .B(n1969), .ZN(n1726) );
  AOI22_X1 U2249 ( .A1(reg4[7]), .A2(n1931), .B1(n1930), .B2(n2830), .ZN(n1993) );
  NOR2_X1 U2246 ( .A1(n1991), .A2(n2843), .ZN(n1980) );
  XNOR2_X1 U2235 ( .A(n1986), .B(n1971), .ZN(n1981) );
  XNOR2_X1 U2223 ( .A(n1981), .B(n1984), .ZN(n1730) );
  NOR2_X1 U2257 ( .A1(reg4[5]), .A2(n1907), .ZN(n1996) );
  NOR2_X1 U2243 ( .A1(n1989), .A2(n1990), .ZN(n1982) );
  AOI222_X1 U2222 ( .A1(p10_muxs_out_2__7_), .A2(n1982), .B1(
        p10_muxs_out_2__7_), .B2(n1983), .C1(n1982), .C2(n1983), .ZN(n1733) );
  XNOR2_X1 U2255 ( .A(p10_muxs_out_1__6_), .B(n1989), .ZN(n1995) );
  NAND2_X1 U2254 ( .A1(n1995), .A2(p10_muxs_out_2__6_), .ZN(n1738) );
  AOI222_X1 U2239 ( .A1(n1736), .A2(n1739), .B1(n1736), .B2(n1738), .C1(n1739), 
        .C2(n1738), .ZN(p10_C[55]) );
  AOI22_X1 U1938 ( .A1(p10_muxs_out_3__7_), .A2(n1737), .B1(n1738), .B2(n1739), 
        .ZN(n1735) );
  XNOR2_X1 U1937 ( .A(n1735), .B(n1736), .ZN(p10_S[55]) );
  OAI21_X1 U2253 ( .B1(n1995), .B2(p10_muxs_out_2__6_), .A(n1738), .ZN(n1740)
         );
  NOR2_X1 U2252 ( .A1(n1994), .A2(n1740), .ZN(p10_C[54]) );
  XNOR2_X1 U1940 ( .A(p10_muxs_out_3__6_), .B(n1740), .ZN(p10_S[54]) );
  AOI222_X1 U2205 ( .A1(n1728), .A2(n1729), .B1(n1728), .B2(n1726), .C1(n1729), 
        .C2(n1726), .ZN(p10_C[57]) );
  AOI22_X1 U1415 ( .A1(reg1_reg[11]), .A2(n2848), .B1(reg1_reg[12]), .B2(n2790), .ZN(n1236) );
  OAI21_X1 U1395 ( .B1(reg1_reg[11]), .B2(reg1_reg[12]), .A(n994), .ZN(n1238)
         );
  AOI22_X1 U1199 ( .A1(B0[12]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_25_), .ZN(n1073) );
  OAI221_X1 U1198 ( .B1(B0[11]), .B2(n993), .C1(n2900), .C2(n994), .A(n1073), 
        .ZN(p6_C[72]) );
  AOI22_X1 U1157 ( .A1(B0[13]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_38_), .ZN(n995) );
  OAI221_X1 U1156 ( .B1(B0[12]), .B2(n993), .C1(p6_minus_A_shifted_25_), .C2(
        n994), .A(n995), .ZN(p6_final_product2_26_) );
  OAI21_X1 U1460 ( .B1(reg1_reg[9]), .B2(reg1_reg[10]), .A(n1075), .ZN(n1274)
         );
  AOI22_X1 U1214 ( .A1(B0[12]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_25_), .ZN(n1092) );
  OAI221_X1 U1213 ( .B1(B0[11]), .B2(n1074), .C1(n2900), .C2(n1075), .A(n1092), 
        .ZN(n1083) );
  OAI21_X1 U1498 ( .B1(reg1_reg[8]), .B2(p6_Partial_products_sum_add_23_B_0_), 
        .A(n1090), .ZN(n1306) );
  AOI22_X1 U1224 ( .A1(B0[13]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_38_), .ZN(n1091) );
  OAI221_X1 U1212 ( .B1(B0[13]), .B2(n1089), .C1(p6_minus_A_shifted_38_), .C2(
        n1090), .A(n1091), .ZN(n1086) );
  AOI22_X1 U1210 ( .A1(B0[10]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_23_), .ZN(n1088) );
  OAI221_X1 U1209 ( .B1(B0[9]), .B2(n993), .C1(p6_minus_A_shifted_22_), .C2(
        n994), .A(n1088), .ZN(n1085) );
  AOI222_X1 U1205 ( .A1(n1083), .A2(n1084), .B1(n1083), .B2(n1085), .C1(n1084), 
        .C2(n1085), .ZN(n1001) );
  AOI22_X1 U1204 ( .A1(B0[11]), .A2(n1081), .B1(n1082), .B2(n2900), .ZN(n1080)
         );
  AOI221_X1 U1203 ( .B1(B0[10]), .B2(n998), .C1(p6_minus_A_shifted_23_), .C2(
        n1079), .A(n1080), .ZN(n1002) );
  AOI22_X1 U1202 ( .A1(B0[13]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_38_), .ZN(n1076) );
  OAI221_X1 U1201 ( .B1(B0[12]), .B2(n1074), .C1(p6_minus_A_shifted_25_), .C2(
        n1075), .A(n1076), .ZN(n999) );
  AOI222_X1 U1200 ( .A1(n1001), .A2(n1002), .B1(n1001), .B2(n999), .C1(n1002), 
        .C2(n999), .ZN(p6_C[71]) );
  XNOR2_X1 U1160 ( .A(n999), .B(n1000), .ZN(p6_S[71]) );
  OAI221_X1 U1223 ( .B1(B0[12]), .B2(n1089), .C1(p6_minus_A_shifted_25_), .C2(
        n1090), .A(n1091), .ZN(n1005) );
  AOI22_X1 U1222 ( .A1(B0[11]), .A2(n1077), .B1(n1078), .B2(n2900), .ZN(n1097)
         );
  OAI221_X1 U1221 ( .B1(B0[10]), .B2(n1074), .C1(p6_minus_A_shifted_23_), .C2(
        n1075), .A(n1097), .ZN(n1093) );
  AOI22_X1 U1245 ( .A1(B0[12]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_25_), .ZN(n1117) );
  OAI221_X1 U1244 ( .B1(B0[11]), .B2(n1089), .C1(n2900), .C2(n1090), .A(n1117), 
        .ZN(n1100) );
  AOI22_X1 U1242 ( .A1(B0[10]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_23_), .ZN(n1116) );
  OAI221_X1 U1241 ( .B1(B0[9]), .B2(n1074), .C1(p6_minus_A_shifted_22_), .C2(
        n1075), .A(n1116), .ZN(n1101) );
  AOI222_X1 U1225 ( .A1(n1100), .A2(n1101), .B1(n1100), .B2(n1102), .C1(n1101), 
        .C2(n1102), .ZN(n1095) );
  AOI222_X1 U1215 ( .A1(n1093), .A2(n1008), .B1(n1093), .B2(n1094), .C1(n1008), 
        .C2(n1094), .ZN(n1004) );
  XNOR2_X1 U1211 ( .A(n1083), .B(n1086), .ZN(n1087) );
  XNOR2_X1 U1208 ( .A(n1087), .B(n1085), .ZN(n1007) );
  AOI222_X1 U1207 ( .A1(n1008), .A2(n1004), .B1(n1008), .B2(n1007), .C1(n1004), 
        .C2(n1007), .ZN(p6_C[70]) );
  AOI22_X1 U1163 ( .A1(n1005), .A2(n1006), .B1(n1007), .B2(n1008), .ZN(n1003)
         );
  XNOR2_X1 U1162 ( .A(n1003), .B(n1004), .ZN(p6_S[70]) );
  XNOR2_X1 U1243 ( .A(p6_muxs_out_3__20_), .B(n1100), .ZN(n1115) );
  AOI22_X1 U1239 ( .A1(B0[8]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_21_), .ZN(n1114) );
  OAI221_X1 U1238 ( .B1(B0[7]), .B2(n993), .C1(p6_minus_A_shifted_20_), .C2(
        n994), .A(n1114), .ZN(n1105) );
  AOI22_X1 U1255 ( .A1(B0[8]), .A2(n1075), .B1(n1074), .B2(
        p6_minus_A_shifted_21_), .ZN(n1124) );
  AOI221_X1 U1254 ( .B1(n1077), .B2(B0[9]), .C1(n1078), .C2(
        p6_minus_A_shifted_22_), .A(n1124), .ZN(n1111) );
  AOI22_X1 U1258 ( .A1(B0[11]), .A2(n1098), .B1(n1099), .B2(n2900), .ZN(n1125)
         );
  OAI221_X1 U1257 ( .B1(B0[10]), .B2(n1089), .C1(p6_minus_A_shifted_23_), .C2(
        n1090), .A(n1125), .ZN(n1113) );
  AOI222_X1 U1235 ( .A1(p6_muxs_out_3__19_), .A2(n1111), .B1(
        p6_muxs_out_3__19_), .B2(n1112), .C1(n1111), .C2(n1112), .ZN(n1106) );
  AOI222_X1 U1229 ( .A1(n1104), .A2(n1105), .B1(n1104), .B2(n1106), .C1(n1105), 
        .C2(n1106), .ZN(n1011) );
  AOI22_X1 U1228 ( .A1(B0[9]), .A2(n1081), .B1(n1082), .B2(
        p6_minus_A_shifted_22_), .ZN(n1103) );
  AOI221_X1 U1227 ( .B1(B0[8]), .B2(n998), .C1(p6_minus_A_shifted_21_), .C2(
        n1079), .A(n1103), .ZN(n1012) );
  XNOR2_X1 U1219 ( .A(n1095), .B(n1096), .ZN(n1009) );
  AOI222_X1 U1218 ( .A1(n1011), .A2(n1012), .B1(n1011), .B2(n1009), .C1(n1012), 
        .C2(n1009), .ZN(p6_C[69]) );
  XNOR2_X1 U1165 ( .A(n1009), .B(n1010), .ZN(p6_S[69]) );
  XNOR2_X1 U1234 ( .A(n1110), .B(n1106), .ZN(n1013) );
  XNOR2_X1 U1256 ( .A(p6_muxs_out_3__19_), .B(n1113), .ZN(n1123) );
  AOI22_X1 U1275 ( .A1(B0[8]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_21_), .ZN(n1138) );
  OAI221_X1 U1274 ( .B1(B0[7]), .B2(n1074), .C1(p6_minus_A_shifted_20_), .C2(
        n1075), .A(n1138), .ZN(n1128) );
  AOI22_X1 U1272 ( .A1(B0[6]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_19_), .ZN(n1137) );
  OAI221_X1 U1271 ( .B1(B0[5]), .B2(n993), .C1(p6_minus_A_shifted_18_), .C2(
        n994), .A(n1137), .ZN(n1129) );
  AOI222_X1 U1263 ( .A1(p6_muxs_out_2__17_), .A2(n1128), .B1(
        p6_muxs_out_2__17_), .B2(n1129), .C1(n1128), .C2(n1129), .ZN(n1108) );
  AOI22_X1 U1279 ( .A1(B0[10]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_23_), .ZN(n1140) );
  OAI221_X1 U1278 ( .B1(B0[9]), .B2(n1089), .C1(p6_minus_A_shifted_22_), .C2(
        n1090), .A(n1140), .ZN(n1126) );
  AOI222_X1 U1261 ( .A1(p6_muxs_out_3__18_), .A2(n1126), .B1(
        p6_muxs_out_3__18_), .B2(n1127), .C1(n1126), .C2(n1127), .ZN(n1109) );
  OAI222_X1 U1232 ( .A1(n1107), .A2(n1108), .B1(n1107), .B2(n1109), .C1(n1108), 
        .C2(n1109), .ZN(n1015) );
  AOI222_X1 U1230 ( .A1(n1013), .A2(n1017), .B1(n1013), .B2(n1016), .C1(n1017), 
        .C2(n1016), .ZN(p6_C[68]) );
  AOI22_X1 U1168 ( .A1(p6_muxs_out_3__19_), .A2(n1015), .B1(n1016), .B2(n1017), 
        .ZN(n1014) );
  XNOR2_X1 U1167 ( .A(n1013), .B(n1014), .ZN(p6_S[68]) );
  XNOR2_X1 U1260 ( .A(n1108), .B(n1109), .ZN(n1122) );
  XNOR2_X1 U1252 ( .A(n1122), .B(n1107), .ZN(n1018) );
  XNOR2_X1 U1273 ( .A(p6_muxs_out_2__17_), .B(n1128), .ZN(n1136) );
  XNOR2_X1 U1270 ( .A(n1136), .B(n1129), .ZN(n1119) );
  AOI222_X1 U1296 ( .A1(p6_muxs_out_2__16_), .A2(p6_muxs_out_3__16_), .B1(
        p6_muxs_out_2__16_), .B2(n1154), .C1(p6_muxs_out_3__16_), .C2(n1154), 
        .ZN(n1135) );
  AOI222_X1 U1268 ( .A1(p6_muxs_out_2__17_), .A2(n1134), .B1(
        p6_muxs_out_2__17_), .B2(n1135), .C1(n1134), .C2(n1135), .ZN(n1120) );
  XNOR2_X1 U1276 ( .A(p6_muxs_out_2__18_), .B(n1139), .ZN(n1121) );
  AOI222_X1 U1251 ( .A1(n1119), .A2(n1120), .B1(n1119), .B2(n1121), .C1(n1120), 
        .C2(n1121), .ZN(n1021) );
  OAI22_X1 U1248 ( .A1(p6_minus_A_shifted_20_), .A2(n1081), .B1(n1082), .B2(
        B0[7]), .ZN(n1118) );
  AOI221_X1 U1247 ( .B1(p6_minus_A_shifted_19_), .B2(n1079), .C1(B0[6]), .C2(
        n998), .A(n1118), .ZN(n1020) );
  AOI222_X1 U1246 ( .A1(n1018), .A2(n1021), .B1(n1018), .B2(n1020), .C1(n1021), 
        .C2(n1020), .ZN(p6_C[67]) );
  XNOR2_X1 U1170 ( .A(n1020), .B(n1021), .ZN(n1019) );
  AOI22_X1 U1293 ( .A1(B0[7]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_20_), .ZN(n1152) );
  OAI221_X1 U1292 ( .B1(B0[6]), .B2(n1074), .C1(p6_minus_A_shifted_19_), .C2(
        n1075), .A(n1152), .ZN(n1130) );
  AOI22_X1 U1291 ( .A1(B0[5]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_18_), .ZN(n1151) );
  OAI221_X1 U1290 ( .B1(B0[4]), .B2(n993), .C1(p6_minus_A_shifted_17_), .C2(
        n994), .A(n1151), .ZN(n1131) );
  AOI22_X1 U1289 ( .A1(B0[9]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_22_), .ZN(n1150) );
  OAI221_X1 U1288 ( .B1(B0[8]), .B2(n1089), .C1(p6_minus_A_shifted_21_), .C2(
        n1090), .A(n1150), .ZN(n1132) );
  XNOR2_X1 U1287 ( .A(n1131), .B(n1132), .ZN(n1149) );
  XNOR2_X1 U1286 ( .A(n1130), .B(n1149), .ZN(n1141) );
  XNOR2_X1 U1307 ( .A(p6_muxs_out_3__16_), .B(p6_muxs_out_2__16_), .ZN(n1163)
         );
  XNOR2_X1 U1306 ( .A(n1163), .B(p6_muxs_out_1__16_), .ZN(n1145) );
  AOI222_X1 U1303 ( .A1(p6_muxs_out_3__15_), .A2(p6_muxs_out_2__15_), .B1(
        p6_muxs_out_3__15_), .B2(n1162), .C1(p6_muxs_out_2__15_), .C2(n1162), 
        .ZN(n1146) );
  AOI22_X1 U1309 ( .A1(B0[8]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_21_), .ZN(n1164) );
  OAI221_X1 U1308 ( .B1(B0[7]), .B2(n1089), .C1(p6_minus_A_shifted_20_), .C2(
        n1090), .A(n1164), .ZN(n1148) );
  AOI222_X1 U1283 ( .A1(n1145), .A2(n1146), .B1(n1145), .B2(n1147), .C1(n1146), 
        .C2(n1147), .ZN(n1143) );
  AOI222_X1 U1280 ( .A1(n1141), .A2(n1142), .B1(n1141), .B2(n1143), .C1(n1142), 
        .C2(n1143), .ZN(n1024) );
  XNOR2_X1 U1266 ( .A(n1121), .B(n1133), .ZN(n1025) );
  AOI222_X1 U1265 ( .A1(n1130), .A2(n1131), .B1(n1130), .B2(n1132), .C1(n1131), 
        .C2(n1132), .ZN(n1022) );
  AOI222_X1 U1264 ( .A1(n1024), .A2(n1025), .B1(n1024), .B2(n1022), .C1(n1025), 
        .C2(n1022), .ZN(p6_C[66]) );
  XNOR2_X1 U1171 ( .A(n1022), .B(n1023), .ZN(p6_S[66]) );
  AOI22_X1 U1317 ( .A1(B0[6]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_19_), .ZN(n1170) );
  OAI221_X1 U1316 ( .B1(B0[5]), .B2(n1074), .C1(p6_minus_A_shifted_18_), .C2(
        n1075), .A(n1170), .ZN(n1158) );
  AOI22_X1 U1315 ( .A1(B0[4]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_17_), .ZN(n1169) );
  OAI221_X1 U1314 ( .B1(B0[3]), .B2(n993), .C1(p6_minus_A_shifted_16_), .C2(
        n994), .A(n1169), .ZN(n1159) );
  AOI222_X1 U1299 ( .A1(p6_muxs_out_1__15_), .A2(n1158), .B1(
        p6_muxs_out_1__15_), .B2(n1159), .C1(n1158), .C2(n1159), .ZN(n1028) );
  XNOR2_X1 U1313 ( .A(n1158), .B(n1159), .ZN(n1168) );
  XNOR2_X1 U1312 ( .A(p6_muxs_out_1__15_), .B(n1168), .ZN(n1155) );
  NOR2_X1 U1529 ( .A1(reg1_reg[1]), .A2(n2836), .ZN(n1212) );
  AOI22_X1 U1357 ( .A1(B0[13]), .A2(n1212), .B1(reg1_reg[1]), .B2(
        p6_minus_A_shifted_38_), .ZN(n1195) );
  NOR2_X1 U1340 ( .A1(p6_muxs_out_1__14_), .A2(n1195), .ZN(n1165) );
  XNOR2_X1 U1339 ( .A(p6_muxs_out_1__15_), .B(p6_muxs_out_3__15_), .ZN(n1194)
         );
  XNOR2_X1 U1338 ( .A(n1194), .B(p6_muxs_out_2__15_), .ZN(n1166) );
  AOI22_X1 U1354 ( .A1(B0[6]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_19_), .ZN(n1211) );
  OAI221_X1 U1353 ( .B1(B0[5]), .B2(n1089), .C1(p6_minus_A_shifted_18_), .C2(
        n1090), .A(n1211), .ZN(n1196) );
  AOI222_X1 U1341 ( .A1(p6_muxs_out_3__14_), .A2(p6_muxs_out_2__14_), .B1(
        p6_muxs_out_3__14_), .B2(n1196), .C1(p6_muxs_out_2__14_), .C2(n1196), 
        .ZN(n1167) );
  AOI222_X1 U1311 ( .A1(n1165), .A2(n1166), .B1(n1165), .B2(n1167), .C1(n1166), 
        .C2(n1167), .ZN(n1156) );
  XNOR2_X1 U1305 ( .A(n1148), .B(n1145), .ZN(n1161) );
  XNOR2_X1 U1302 ( .A(n1161), .B(n1146), .ZN(n1157) );
  AOI222_X1 U1298 ( .A1(n1155), .A2(n1156), .B1(n1155), .B2(n1157), .C1(n1156), 
        .C2(n1157), .ZN(n1029) );
  XNOR2_X1 U1282 ( .A(n1144), .B(n1143), .ZN(n1026) );
  AOI222_X1 U1281 ( .A1(n1028), .A2(n1029), .B1(n1028), .B2(n1026), .C1(n1029), 
        .C2(n1026), .ZN(p6_C[65]) );
  XNOR2_X1 U1173 ( .A(n1026), .B(n1027), .ZN(p6_S[65]) );
  AOI22_X1 U1335 ( .A1(B0[5]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_18_), .ZN(n1192) );
  OAI221_X1 U1334 ( .B1(B0[4]), .B2(n1074), .C1(p6_minus_A_shifted_17_), .C2(
        n1075), .A(n1192), .ZN(n1174) );
  AOI22_X1 U1333 ( .A1(B0[3]), .A2(n996), .B1(n997), .B2(
        p6_minus_A_shifted_16_), .ZN(n1191) );
  OAI221_X1 U1332 ( .B1(B0[2]), .B2(n993), .C1(p6_minus_A_shifted_15_), .C2(
        n994), .A(n1191), .ZN(n1175) );
  AOI22_X1 U1330 ( .A1(B0[7]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_20_), .ZN(n1190) );
  OAI221_X1 U1329 ( .B1(B0[6]), .B2(n1089), .C1(p6_minus_A_shifted_19_), .C2(
        n1090), .A(n1190), .ZN(n1176) );
  AOI222_X1 U1319 ( .A1(n1174), .A2(n1175), .B1(n1174), .B2(n1176), .C1(n1175), 
        .C2(n1176), .ZN(n1032) );
  XNOR2_X1 U1331 ( .A(n1174), .B(n1175), .ZN(n1189) );
  XNOR2_X1 U1328 ( .A(n1189), .B(n1176), .ZN(n1171) );
  XNOR2_X1 U1336 ( .A(n1167), .B(n1193), .ZN(n1172) );
  NAND2_X1 U1525 ( .A1(reg1_reg[1]), .A2(n2836), .ZN(n1228) );
  NAND2_X1 U1527 ( .A1(reg1_reg[0]), .A2(reg1_reg[1]), .ZN(n1246) );
  AOI22_X1 U1379 ( .A1(B0[13]), .A2(n1212), .B1(n1230), .B2(
        p6_minus_A_shifted_38_), .ZN(n1229) );
  OAI21_X1 U1378 ( .B1(B0[12]), .B2(n1228), .A(n1229), .ZN(n1227) );
  NAND2_X1 U1377 ( .A1(n1227), .A2(p6_muxs_out_1__13_), .ZN(n1186) );
  XNOR2_X1 U1355 ( .A(p6_muxs_out_3__14_), .B(p6_muxs_out_2__14_), .ZN(n1210)
         );
  OAI222_X1 U1326 ( .A1(n1186), .A2(n1187), .B1(n1186), .B2(n1188), .C1(n1187), 
        .C2(n1188), .ZN(n1173) );
  AOI222_X1 U1318 ( .A1(n1171), .A2(n1172), .B1(n1171), .B2(n1173), .C1(n1172), 
        .C2(n1173), .ZN(n1031) );
  XNOR2_X1 U1310 ( .A(n1155), .B(n1156), .ZN(n1160) );
  AOI222_X1 U1300 ( .A1(n1032), .A2(n1031), .B1(n1032), .B2(n1033), .C1(n1031), 
        .C2(n1033), .ZN(p6_C[64]) );
  XNOR2_X1 U1175 ( .A(n1030), .B(n1031), .ZN(p6_S[64]) );
  XNOR2_X1 U1327 ( .A(n1172), .B(n1171), .ZN(n1185) );
  XNOR2_X1 U1351 ( .A(n1187), .B(n1188), .ZN(n1209) );
  AOI22_X1 U1384 ( .A1(B0[5]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_18_), .ZN(n1232) );
  OAI221_X1 U1383 ( .B1(B0[4]), .B2(n1089), .C1(p6_minus_A_shifted_17_), .C2(
        n1090), .A(n1232), .ZN(n1216) );
  AOI222_X1 U1364 ( .A1(p6_muxs_out_2__13_), .A2(p6_muxs_out_3__13_), .B1(
        p6_muxs_out_2__13_), .B2(n1216), .C1(p6_muxs_out_3__13_), .C2(n1216), 
        .ZN(n1179) );
  AOI22_X1 U1363 ( .A1(B0[1]), .A2(n994), .B1(n993), .B2(
        p6_minus_A_shifted_14_), .ZN(n1215) );
  AOI221_X1 U1362 ( .B1(n996), .B2(B0[2]), .C1(n997), .C2(
        p6_minus_A_shifted_15_), .A(n1215), .ZN(n1180) );
  XNOR2_X1 U1361 ( .A(n1179), .B(n1180), .ZN(n1213) );
  AOI22_X1 U1360 ( .A1(B0[4]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_17_), .ZN(n1214) );
  OAI221_X1 U1359 ( .B1(B0[3]), .B2(n1074), .C1(p6_minus_A_shifted_16_), .C2(
        n1075), .A(n1214), .ZN(n1181) );
  XNOR2_X1 U1358 ( .A(n1213), .B(n1181), .ZN(n1183) );
  XNOR2_X1 U1381 ( .A(p6_muxs_out_2__13_), .B(n1231), .ZN(n1206) );
  OAI21_X1 U1376 ( .B1(n1227), .B2(p6_muxs_out_1__13_), .A(n1186), .ZN(n1207)
         );
  OAI222_X1 U1406 ( .A1(B0[12]), .A2(n1246), .B1(p6_minus_A_shifted_25_), .B2(
        n1247), .C1(B0[11]), .C2(n1228), .ZN(n1245) );
  NAND2_X1 U1405 ( .A1(n1245), .A2(p6_muxs_out_1__12_), .ZN(n1208) );
  AOI222_X1 U1348 ( .A1(n1206), .A2(n1207), .B1(n1206), .B2(n1208), .C1(n1207), 
        .C2(n1208), .ZN(n1184) );
  AOI222_X1 U1324 ( .A1(n1182), .A2(n1183), .B1(n1182), .B2(n1184), .C1(n1183), 
        .C2(n1184), .ZN(n1037) );
  OAI222_X1 U1322 ( .A1(n1178), .A2(n1179), .B1(n1178), .B2(n1180), .C1(n1179), 
        .C2(n1180), .ZN(n1177) );
  AOI222_X1 U1320 ( .A1(n1036), .A2(n1037), .B1(n1036), .B2(n1034), .C1(n1037), 
        .C2(n1034), .ZN(p6_C[63]) );
  XNOR2_X1 U1177 ( .A(n1034), .B(n1035), .ZN(p6_S[63]) );
  XNOR2_X1 U1347 ( .A(n1205), .B(n1184), .ZN(n1040) );
  XNOR2_X1 U1375 ( .A(n1206), .B(n1207), .ZN(n1226) );
  AOI22_X1 U1411 ( .A1(B0[4]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_17_), .ZN(n1249) );
  OAI221_X1 U1410 ( .B1(B0[3]), .B2(n1089), .C1(p6_minus_A_shifted_16_), .C2(
        n1090), .A(n1249), .ZN(n1239) );
  AOI222_X1 U1397 ( .A1(p6_muxs_out_2__12_), .A2(p6_muxs_out_3__12_), .B1(
        p6_muxs_out_2__12_), .B2(n1239), .C1(p6_muxs_out_3__12_), .C2(n1239), 
        .ZN(n1199) );
  AOI22_X1 U1391 ( .A1(B0[0]), .A2(n994), .B1(n993), .B2(
        p6_minus_A_shifted_13_), .ZN(n1235) );
  AOI221_X1 U1390 ( .B1(n996), .B2(B0[1]), .C1(n997), .C2(
        p6_minus_A_shifted_14_), .A(n1235), .ZN(n1200) );
  XNOR2_X1 U1389 ( .A(n1199), .B(n1200), .ZN(n1233) );
  AOI22_X1 U1388 ( .A1(B0[3]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_16_), .ZN(n1234) );
  OAI221_X1 U1387 ( .B1(B0[2]), .B2(n1074), .C1(p6_minus_A_shifted_15_), .C2(
        n1075), .A(n1234), .ZN(n1201) );
  XNOR2_X1 U1386 ( .A(n1233), .B(n1201), .ZN(n1203) );
  XNOR2_X1 U1408 ( .A(p6_muxs_out_2__12_), .B(n1248), .ZN(n1223) );
  OAI21_X1 U1404 ( .B1(n1245), .B2(p6_muxs_out_1__12_), .A(n1208), .ZN(n1224)
         );
  AOI22_X1 U1430 ( .A1(n1269), .A2(p6_minus_A_shifted_23_), .B1(n1212), .B2(
        B0[11]), .ZN(n1268) );
  OAI21_X1 U1429 ( .B1(B0[11]), .B2(n1246), .A(n1268), .ZN(n1267) );
  NAND2_X1 U1428 ( .A1(p6_muxs_out_1__11_), .A2(n1267), .ZN(n1225) );
  AOI222_X1 U1372 ( .A1(n1223), .A2(n1224), .B1(n1223), .B2(n1225), .C1(n1224), 
        .C2(n1225), .ZN(n1204) );
  AOI222_X1 U1346 ( .A1(n1202), .A2(n1203), .B1(n1202), .B2(n1204), .C1(n1203), 
        .C2(n1204), .ZN(n1041) );
  OAI222_X1 U1344 ( .A1(n1198), .A2(n1199), .B1(n1198), .B2(n1200), .C1(n1199), 
        .C2(n1200), .ZN(n1197) );
  AOI222_X1 U1342 ( .A1(n1040), .A2(n1041), .B1(n1040), .B2(n1038), .C1(n1041), 
        .C2(n1038), .ZN(p6_C[62]) );
  XNOR2_X1 U1179 ( .A(n1038), .B(n1039), .ZN(p6_S[62]) );
  XNOR2_X1 U1371 ( .A(n1222), .B(n1204), .ZN(n1044) );
  AOI22_X1 U1417 ( .A1(B0[2]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_15_), .ZN(n1253) );
  OAI221_X1 U1416 ( .B1(B0[1]), .B2(n1074), .C1(p6_minus_A_shifted_14_), .C2(
        n1075), .A(n1253), .ZN(n1217) );
  NOR2_X1 U1414 ( .A1(n1236), .A2(p6_minus_A_shifted_13_), .ZN(n1250) );
  XNOR2_X1 U1403 ( .A(n1223), .B(n1224), .ZN(n1244) );
  OAI21_X1 U1427 ( .B1(p6_muxs_out_1__11_), .B2(n1267), .A(n1225), .ZN(n1254)
         );
  AOI22_X1 U1454 ( .A1(n1269), .A2(p6_minus_A_shifted_22_), .B1(n1212), .B2(
        B0[10]), .ZN(n1282) );
  OAI21_X1 U1453 ( .B1(B0[10]), .B2(n1246), .A(n1282), .ZN(n1281) );
  NAND2_X1 U1452 ( .A1(p6_muxs_out_1__10_), .A2(n1281), .ZN(n1256) );
  AOI222_X1 U1418 ( .A1(n1254), .A2(n1255), .B1(n1254), .B2(n1256), .C1(n1255), 
        .C2(n1256), .ZN(n1221) );
  AOI222_X1 U1370 ( .A1(n1219), .A2(n1220), .B1(n1219), .B2(n1221), .C1(n1220), 
        .C2(n1221), .ZN(n1045) );
  OAI221_X1 U1367 ( .B1(B0[0]), .B2(n1082), .C1(p6_minus_A_shifted_13_), .C2(
        n1081), .A(n993), .ZN(n1218) );
  AOI222_X1 U1366 ( .A1(n1217), .A2(reg1_reg[13]), .B1(n1217), .B2(n1218), 
        .C1(reg1_reg[13]), .C2(n1218), .ZN(n1042) );
  AOI222_X1 U1365 ( .A1(n1044), .A2(n1045), .B1(n1044), .B2(n1042), .C1(n1045), 
        .C2(n1042), .ZN(p6_C[61]) );
  XNOR2_X1 U1181 ( .A(n1042), .B(n1043), .ZN(p6_S[61]) );
  AOI22_X1 U1441 ( .A1(B0[1]), .A2(n1077), .B1(n1078), .B2(
        p6_minus_A_shifted_14_), .ZN(n1273) );
  OAI221_X1 U1440 ( .B1(B0[0]), .B2(n1074), .C1(p6_minus_A_shifted_13_), .C2(
        n1075), .A(n1273), .ZN(n1257) );
  AOI22_X1 U1437 ( .A1(B0[3]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_16_), .ZN(n1272) );
  OAI221_X1 U1436 ( .B1(B0[2]), .B2(n1089), .C1(p6_minus_A_shifted_15_), .C2(
        n1090), .A(n1272), .ZN(n1258) );
  AOI222_X1 U1419 ( .A1(n1257), .A2(p6_muxs_out_3__11_), .B1(n1257), .B2(n1258), .C1(p6_muxs_out_3__11_), .C2(n1258), .ZN(n1048) );
  XNOR2_X1 U1400 ( .A(n1221), .B(n1243), .ZN(n1049) );
  XNOR2_X1 U1439 ( .A(n1257), .B(p6_muxs_out_3__11_), .ZN(n1271) );
  XNOR2_X1 U1435 ( .A(n1271), .B(n1258), .ZN(n1240) );
  AOI22_X1 U1432 ( .A1(p6_muxs_out_2__11_), .A2(n1270), .B1(n1256), .B2(n1255), 
        .ZN(n1266) );
  XNOR2_X1 U1426 ( .A(n1266), .B(n1254), .ZN(n1241) );
  OAI21_X1 U1451 ( .B1(p6_muxs_out_1__10_), .B2(n1281), .A(n1256), .ZN(n1277)
         );
  AOI222_X1 U1445 ( .A1(n1275), .A2(n1276), .B1(n1275), .B2(n1277), .C1(n1276), 
        .C2(n1277), .ZN(n1242) );
  AOI222_X1 U1399 ( .A1(n1240), .A2(n1241), .B1(n1240), .B2(n1242), .C1(n1241), 
        .C2(n1242), .ZN(n1046) );
  AOI222_X1 U1398 ( .A1(n1048), .A2(n1049), .B1(n1048), .B2(n1046), .C1(n1049), 
        .C2(n1046), .ZN(p6_C[60]) );
  AOI22_X1 U1481 ( .A1(p6_muxs_out_1__9_), .A2(p6_muxs_out_2__9_), .B1(n1285), 
        .B2(n1284), .ZN(n1297) );
  NOR2_X1 U1479 ( .A1(B0[8]), .A2(n1228), .ZN(n1298) );
  AOI221_X1 U1478 ( .B1(B0[9]), .B2(n1212), .C1(p6_minus_A_shifted_22_), .C2(
        n1230), .A(n1298), .ZN(n1286) );
  XNOR2_X1 U1477 ( .A(n1297), .B(n1286), .ZN(n1287) );
  AOI22_X1 U1475 ( .A1(B0[0]), .A2(n1090), .B1(n1089), .B2(
        p6_minus_A_shifted_13_), .ZN(n1296) );
  OAI221_X1 U1473 ( .B1(n1293), .B2(p6_minus_A_shifted_14_), .C1(n1294), .C2(
        B0[1]), .A(n1295), .ZN(n1278) );
  AOI22_X1 U1502 ( .A1(B0[8]), .A2(n1212), .B1(n1230), .B2(
        p6_minus_A_shifted_21_), .ZN(n1308) );
  OAI21_X1 U1501 ( .B1(B0[7]), .B2(n1228), .A(n1308), .ZN(n1292) );
  AOI222_X1 U1470 ( .A1(p6_muxs_out_1__8_), .A2(p6_muxs_out_2__8_), .B1(
        p6_muxs_out_1__8_), .B2(n1292), .C1(p6_muxs_out_2__8_), .C2(n1292), 
        .ZN(n1290) );
  AOI222_X1 U1466 ( .A1(n1287), .A2(n1288), .B1(n1287), .B2(n1289), .C1(n1288), 
        .C2(n1289), .ZN(n1056) );
  AOI222_X1 U1465 ( .A1(n1284), .A2(n1285), .B1(n1284), .B2(n1286), .C1(n1285), 
        .C2(n1286), .ZN(n1264) );
  AOI22_X1 U1463 ( .A1(B0[2]), .A2(n1098), .B1(n1099), .B2(
        p6_minus_A_shifted_15_), .ZN(n1283) );
  OAI221_X1 U1462 ( .B1(B0[1]), .B2(n1089), .C1(p6_minus_A_shifted_14_), .C2(
        n1090), .A(n1283), .ZN(n1260) );
  NOR2_X1 U1459 ( .A1(n1274), .A2(p6_minus_A_shifted_13_), .ZN(n1261) );
  AOI22_X1 U1455 ( .A1(p6_muxs_out_2__10_), .A2(p6_muxs_out_3__10_), .B1(n1276), .B2(n1275), .ZN(n1280) );
  XNOR2_X1 U1450 ( .A(n1280), .B(n1277), .ZN(n1263) );
  XNOR2_X1 U1448 ( .A(n1264), .B(n1279), .ZN(n1057) );
  NAND2_X1 U1447 ( .A1(p6_muxs_out_3__9_), .A2(n1278), .ZN(n1054) );
  AOI222_X1 U1446 ( .A1(n1056), .A2(n1057), .B1(n1056), .B2(n1054), .C1(n1057), 
        .C2(n1054), .ZN(p6_C[58]) );
  XNOR2_X1 U1424 ( .A(n1242), .B(n1265), .ZN(n1052) );
  AOI222_X1 U1423 ( .A1(n1262), .A2(n1263), .B1(n1262), .B2(n1264), .C1(n1263), 
        .C2(n1264), .ZN(n1053) );
  XNOR2_X1 U1185 ( .A(n1050), .B(n1051), .ZN(p6_S[59]) );
  XNOR2_X1 U1504 ( .A(p6_muxs_out_2__8_), .B(p6_muxs_out_1__8_), .ZN(n1307) );
  XNOR2_X1 U1500 ( .A(n1307), .B(n1292), .ZN(n1302) );
  OAI221_X1 U1491 ( .B1(n1293), .B2(p6_minus_A_shifted_13_), .C1(n1294), .C2(
        B0[0]), .A(n1089), .ZN(n1299) );
  AOI22_X1 U1515 ( .A1(B0[7]), .A2(n1247), .B1(n1246), .B2(
        p6_minus_A_shifted_20_), .ZN(n1314) );
  AOI21_X1 U1514 ( .B1(n1269), .B2(p6_minus_A_shifted_19_), .A(n1314), .ZN(
        n1312) );
  NOR2_X1 U1512 ( .A1(n1312), .A2(n2850), .ZN(n1301) );
  XNOR2_X1 U1488 ( .A(n1302), .B(n1305), .ZN(n1062) );
  NOR2_X1 U1524 ( .A1(B0[5]), .A2(n1228), .ZN(n1317) );
  AOI221_X1 U1523 ( .B1(B0[6]), .B2(n1212), .C1(p6_minus_A_shifted_19_), .C2(
        n1230), .A(n1317), .ZN(n1310) );
  NOR2_X1 U1509 ( .A1(n1310), .A2(n1311), .ZN(n1303) );
  AOI21_X1 U1511 ( .B1(n1312), .B2(n2850), .A(n1301), .ZN(n1304) );
  AOI222_X1 U1487 ( .A1(p6_muxs_out_2__7_), .A2(n1303), .B1(p6_muxs_out_2__7_), 
        .B2(n1304), .C1(n1303), .C2(n1304), .ZN(n1065) );
  XNOR2_X1 U1471 ( .A(n1287), .B(n1288), .ZN(n1291) );
  XNOR2_X1 U1469 ( .A(n1291), .B(n1290), .ZN(n1058) );
  AOI222_X1 U1485 ( .A1(n1300), .A2(n1301), .B1(n1300), .B2(n1302), .C1(n1301), 
        .C2(n1302), .ZN(n1060) );
  NAND2_X1 U1484 ( .A1(p6_muxs_out_3__8_), .A2(n1299), .ZN(n1061) );
  XNOR2_X1 U1189 ( .A(n1058), .B(n1059), .ZN(p6_S[57]) );
  XNOR2_X1 U1522 ( .A(p6_muxs_out_1__6_), .B(n1310), .ZN(n1316) );
  NAND2_X1 U1521 ( .A1(n1316), .A2(p6_muxs_out_2__6_), .ZN(n1070) );
  OAI21_X1 U1520 ( .B1(n1316), .B2(p6_muxs_out_2__6_), .A(n1070), .ZN(n1072)
         );
  NOR2_X1 U1519 ( .A1(n1315), .A2(n1072), .ZN(p6_C[54]) );
  AOI22_X1 U1195 ( .A1(p6_muxs_out_3__7_), .A2(n1069), .B1(n1070), .B2(n1071), 
        .ZN(n1067) );
  XNOR2_X1 U1507 ( .A(n1304), .B(n1309), .ZN(n1068) );
  XNOR2_X1 U1194 ( .A(n1067), .B(n1068), .ZN(p6_S[55]) );
  XNOR2_X1 U1197 ( .A(p6_muxs_out_3__6_), .B(n1072), .ZN(p6_S[54]) );
  XNOR2_X1 U1191 ( .A(n1062), .B(n1063), .ZN(p6_S[56]) );
  AOI222_X1 U1505 ( .A1(n1068), .A2(n1071), .B1(n1068), .B2(n1070), .C1(n1071), 
        .C2(n1070), .ZN(p6_C[55]) );
  XNOR2_X1 U1187 ( .A(n1054), .B(n1055), .ZN(p6_S[58]) );
  AOI222_X1 U1468 ( .A1(n1060), .A2(n1061), .B1(n1060), .B2(n1058), .C1(n1061), 
        .C2(n1058), .ZN(p6_C[57]) );
  XNOR2_X1 U1183 ( .A(n1046), .B(n1047), .ZN(p6_S[60]) );
  AOI222_X1 U1420 ( .A1(n1052), .A2(n1053), .B1(n1052), .B2(n1050), .C1(n1053), 
        .C2(n1050), .ZN(p6_C[59]) );
  OAI21_X1 U643 ( .B1(reg3_reg[11]), .B2(reg3_reg[12]), .A(n342), .ZN(n586) );
  AOI22_X1 U663 ( .A1(reg3_reg[11]), .A2(n2802), .B1(reg3_reg[12]), .B2(n2786), 
        .ZN(n584) );
  AOI22_X1 U405 ( .A1(B2[13]), .A2(n344), .B1(n345), .B2(
        p8_minus_A_shifted_38_), .ZN(n343) );
  OAI221_X1 U404 ( .B1(B2[12]), .B2(n341), .C1(p8_minus_A_shifted_25_), .C2(
        n342), .A(n343), .ZN(p8_final_product2_26_) );
  AOI22_X1 U447 ( .A1(B2[12]), .A2(n344), .B1(n345), .B2(
        p8_minus_A_shifted_25_), .ZN(n421) );
  OAI221_X1 U446 ( .B1(B2[11]), .B2(n341), .C1(n3068), .C2(n342), .A(n421), 
        .ZN(p8_C[72]) );
  OAI21_X1 U708 ( .B1(reg3_reg[9]), .B2(reg3_reg[10]), .A(n423), .ZN(n622) );
  AOI22_X1 U462 ( .A1(B2[12]), .A2(n425), .B1(n426), .B2(
        p8_minus_A_shifted_25_), .ZN(n440) );
  OAI221_X1 U461 ( .B1(B2[11]), .B2(n422), .C1(n3068), .C2(n423), .A(n440), 
        .ZN(n431) );
  OAI21_X1 U746 ( .B1(reg3_reg[8]), .B2(p8_Partial_products_sum_add_23_B_0_), 
        .A(n438), .ZN(n654) );
  AOI22_X1 U472 ( .A1(B2[13]), .A2(n446), .B1(n447), .B2(
        p8_minus_A_shifted_38_), .ZN(n439) );
  OAI221_X1 U460 ( .B1(B2[13]), .B2(n437), .C1(p8_minus_A_shifted_38_), .C2(
        n438), .A(n439), .ZN(n434) );
  AOI22_X1 U458 ( .A1(B2[10]), .A2(n344), .B1(n345), .B2(
        p8_minus_A_shifted_23_), .ZN(n436) );
  OAI221_X1 U457 ( .B1(B2[9]), .B2(n341), .C1(p8_minus_A_shifted_22_), .C2(
        n342), .A(n436), .ZN(n433) );
  AOI222_X1 U453 ( .A1(n431), .A2(n432), .B1(n431), .B2(n433), .C1(n432), .C2(
        n433), .ZN(n349) );
  AOI22_X1 U452 ( .A1(B2[11]), .A2(n429), .B1(n430), .B2(n3068), .ZN(n428) );
  AOI221_X1 U451 ( .B1(B2[10]), .B2(n346), .C1(p8_minus_A_shifted_23_), .C2(
        n427), .A(n428), .ZN(n350) );
  AOI22_X1 U450 ( .A1(B2[13]), .A2(n425), .B1(n426), .B2(
        p8_minus_A_shifted_38_), .ZN(n424) );
  OAI221_X1 U449 ( .B1(B2[12]), .B2(n422), .C1(p8_minus_A_shifted_25_), .C2(
        n423), .A(n424), .ZN(n347) );
  AOI222_X1 U448 ( .A1(n349), .A2(n350), .B1(n349), .B2(n347), .C1(n350), .C2(
        n347), .ZN(p8_C[71]) );
  XNOR2_X1 U408 ( .A(n347), .B(n348), .ZN(p8_S[71]) );
  OAI221_X1 U471 ( .B1(B2[12]), .B2(n437), .C1(p8_minus_A_shifted_25_), .C2(
        n438), .A(n439), .ZN(n353) );
  AOI22_X1 U470 ( .A1(B2[11]), .A2(n425), .B1(n426), .B2(n3068), .ZN(n445) );
  OAI221_X1 U469 ( .B1(B2[10]), .B2(n422), .C1(p8_minus_A_shifted_23_), .C2(
        n423), .A(n445), .ZN(n441) );
  AOI22_X1 U493 ( .A1(B2[12]), .A2(n446), .B1(n447), .B2(
        p8_minus_A_shifted_25_), .ZN(n465) );
  OAI221_X1 U492 ( .B1(B2[11]), .B2(n437), .C1(n3068), .C2(n438), .A(n465), 
        .ZN(n448) );
  AOI22_X1 U490 ( .A1(B2[10]), .A2(n425), .B1(n426), .B2(
        p8_minus_A_shifted_23_), .ZN(n464) );
  OAI221_X1 U489 ( .B1(B2[9]), .B2(n422), .C1(p8_minus_A_shifted_22_), .C2(
        n423), .A(n464), .ZN(n449) );
  AOI222_X1 U473 ( .A1(n448), .A2(n449), .B1(n448), .B2(n450), .C1(n449), .C2(
        n450), .ZN(n443) );
  AOI222_X1 U463 ( .A1(n441), .A2(n356), .B1(n441), .B2(n442), .C1(n356), .C2(
        n442), .ZN(n352) );
  XNOR2_X1 U459 ( .A(n431), .B(n434), .ZN(n435) );
  XNOR2_X1 U456 ( .A(n435), .B(n433), .ZN(n355) );
  AOI222_X1 U455 ( .A1(n356), .A2(n352), .B1(n356), .B2(n355), .C1(n352), .C2(
        n355), .ZN(p8_C[70]) );
  AOI22_X1 U411 ( .A1(n353), .A2(n354), .B1(n355), .B2(n356), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n351), .B(n352), .ZN(p8_S[70]) );
  XNOR2_X1 U491 ( .A(p8_muxs_out_3__20_), .B(n448), .ZN(n463) );
  AOI22_X1 U487 ( .A1(B2[8]), .A2(n344), .B1(n345), .B2(p8_minus_A_shifted_21_), .ZN(n462) );
  OAI221_X1 U486 ( .B1(B2[7]), .B2(n341), .C1(p8_minus_A_shifted_20_), .C2(
        n342), .A(n462), .ZN(n453) );
  AOI22_X1 U503 ( .A1(B2[8]), .A2(n423), .B1(n422), .B2(p8_minus_A_shifted_21_), .ZN(n472) );
  AOI221_X1 U502 ( .B1(n425), .B2(B2[9]), .C1(n426), .C2(
        p8_minus_A_shifted_22_), .A(n472), .ZN(n459) );
  AOI22_X1 U506 ( .A1(B2[11]), .A2(n446), .B1(n447), .B2(n3068), .ZN(n473) );
  OAI221_X1 U505 ( .B1(B2[10]), .B2(n437), .C1(p8_minus_A_shifted_23_), .C2(
        n438), .A(n473), .ZN(n461) );
  AOI222_X1 U483 ( .A1(p8_muxs_out_3__19_), .A2(n459), .B1(p8_muxs_out_3__19_), 
        .B2(n460), .C1(n459), .C2(n460), .ZN(n454) );
  AOI222_X1 U477 ( .A1(n452), .A2(n453), .B1(n452), .B2(n454), .C1(n453), .C2(
        n454), .ZN(n359) );
  AOI22_X1 U476 ( .A1(B2[9]), .A2(n429), .B1(n430), .B2(p8_minus_A_shifted_22_), .ZN(n451) );
  AOI221_X1 U475 ( .B1(B2[8]), .B2(n346), .C1(p8_minus_A_shifted_21_), .C2(
        n427), .A(n451), .ZN(n360) );
  XNOR2_X1 U467 ( .A(n443), .B(n444), .ZN(n357) );
  AOI222_X1 U466 ( .A1(n359), .A2(n360), .B1(n359), .B2(n357), .C1(n360), .C2(
        n357), .ZN(p8_C[69]) );
  XNOR2_X1 U413 ( .A(n357), .B(n358), .ZN(p8_S[69]) );
  XNOR2_X1 U482 ( .A(n458), .B(n454), .ZN(n361) );
  XNOR2_X1 U504 ( .A(p8_muxs_out_3__19_), .B(n461), .ZN(n471) );
  AOI22_X1 U523 ( .A1(B2[8]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_21_), .ZN(n486) );
  OAI221_X1 U522 ( .B1(B2[7]), .B2(n422), .C1(p8_minus_A_shifted_20_), .C2(
        n423), .A(n486), .ZN(n476) );
  AOI22_X1 U520 ( .A1(B2[6]), .A2(n344), .B1(n345), .B2(p8_minus_A_shifted_19_), .ZN(n485) );
  OAI221_X1 U519 ( .B1(B2[5]), .B2(n341), .C1(p8_minus_A_shifted_18_), .C2(
        n342), .A(n485), .ZN(n477) );
  AOI222_X1 U511 ( .A1(p8_muxs_out_2__17_), .A2(n476), .B1(p8_muxs_out_2__17_), 
        .B2(n477), .C1(n476), .C2(n477), .ZN(n456) );
  AOI22_X1 U527 ( .A1(B2[10]), .A2(n446), .B1(n447), .B2(
        p8_minus_A_shifted_23_), .ZN(n488) );
  OAI221_X1 U526 ( .B1(B2[9]), .B2(n437), .C1(p8_minus_A_shifted_22_), .C2(
        n438), .A(n488), .ZN(n474) );
  AOI222_X1 U509 ( .A1(p8_muxs_out_3__18_), .A2(n474), .B1(p8_muxs_out_3__18_), 
        .B2(n475), .C1(n474), .C2(n475), .ZN(n457) );
  OAI222_X1 U480 ( .A1(n455), .A2(n456), .B1(n455), .B2(n457), .C1(n456), .C2(
        n457), .ZN(n363) );
  AOI222_X1 U478 ( .A1(n361), .A2(n365), .B1(n361), .B2(n364), .C1(n365), .C2(
        n364), .ZN(p8_C[68]) );
  AOI22_X1 U416 ( .A1(p8_muxs_out_3__19_), .A2(n363), .B1(n364), .B2(n365), 
        .ZN(n362) );
  XNOR2_X1 U415 ( .A(n361), .B(n362), .ZN(p8_S[68]) );
  XNOR2_X1 U508 ( .A(n456), .B(n457), .ZN(n470) );
  XNOR2_X1 U500 ( .A(n470), .B(n455), .ZN(n366) );
  XNOR2_X1 U521 ( .A(p8_muxs_out_2__17_), .B(n476), .ZN(n484) );
  XNOR2_X1 U518 ( .A(n484), .B(n477), .ZN(n467) );
  AOI222_X1 U544 ( .A1(p8_muxs_out_2__16_), .A2(p8_muxs_out_3__16_), .B1(
        p8_muxs_out_2__16_), .B2(n502), .C1(p8_muxs_out_3__16_), .C2(n502), 
        .ZN(n483) );
  AOI222_X1 U516 ( .A1(p8_muxs_out_2__17_), .A2(n482), .B1(p8_muxs_out_2__17_), 
        .B2(n483), .C1(n482), .C2(n483), .ZN(n468) );
  XNOR2_X1 U524 ( .A(p8_muxs_out_2__18_), .B(n487), .ZN(n469) );
  AOI222_X1 U499 ( .A1(n467), .A2(n468), .B1(n467), .B2(n469), .C1(n468), .C2(
        n469), .ZN(n369) );
  OAI22_X1 U496 ( .A1(p8_minus_A_shifted_20_), .A2(n429), .B1(n430), .B2(B2[7]), .ZN(n466) );
  AOI221_X1 U495 ( .B1(p8_minus_A_shifted_19_), .B2(n427), .C1(B2[6]), .C2(
        n346), .A(n466), .ZN(n368) );
  AOI222_X1 U494 ( .A1(n366), .A2(n369), .B1(n366), .B2(n368), .C1(n369), .C2(
        n368), .ZN(p8_C[67]) );
  XNOR2_X1 U418 ( .A(n368), .B(n369), .ZN(n367) );
  AOI22_X1 U541 ( .A1(B2[7]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_20_), .ZN(n500) );
  OAI221_X1 U540 ( .B1(B2[6]), .B2(n422), .C1(p8_minus_A_shifted_19_), .C2(
        n423), .A(n500), .ZN(n478) );
  AOI22_X1 U539 ( .A1(B2[5]), .A2(n344), .B1(n345), .B2(p8_minus_A_shifted_18_), .ZN(n499) );
  OAI221_X1 U538 ( .B1(B2[4]), .B2(n341), .C1(p8_minus_A_shifted_17_), .C2(
        n342), .A(n499), .ZN(n479) );
  AOI22_X1 U537 ( .A1(B2[9]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_22_), .ZN(n498) );
  OAI221_X1 U536 ( .B1(B2[8]), .B2(n437), .C1(p8_minus_A_shifted_21_), .C2(
        n438), .A(n498), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n479), .B(n480), .ZN(n497) );
  XNOR2_X1 U534 ( .A(n478), .B(n497), .ZN(n489) );
  XNOR2_X1 U555 ( .A(p8_muxs_out_3__16_), .B(p8_muxs_out_2__16_), .ZN(n511) );
  XNOR2_X1 U554 ( .A(n511), .B(p8_muxs_out_1__16_), .ZN(n493) );
  AOI222_X1 U551 ( .A1(p8_muxs_out_3__15_), .A2(p8_muxs_out_2__15_), .B1(
        p8_muxs_out_3__15_), .B2(n510), .C1(p8_muxs_out_2__15_), .C2(n510), 
        .ZN(n494) );
  AOI22_X1 U557 ( .A1(B2[8]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_21_), .ZN(n512) );
  OAI221_X1 U556 ( .B1(B2[7]), .B2(n437), .C1(p8_minus_A_shifted_20_), .C2(
        n438), .A(n512), .ZN(n496) );
  AOI222_X1 U531 ( .A1(n493), .A2(n494), .B1(n493), .B2(n495), .C1(n494), .C2(
        n495), .ZN(n491) );
  AOI222_X1 U528 ( .A1(n489), .A2(n490), .B1(n489), .B2(n491), .C1(n490), .C2(
        n491), .ZN(n372) );
  XNOR2_X1 U514 ( .A(n469), .B(n481), .ZN(n373) );
  AOI222_X1 U513 ( .A1(n478), .A2(n479), .B1(n478), .B2(n480), .C1(n479), .C2(
        n480), .ZN(n370) );
  AOI222_X1 U512 ( .A1(n372), .A2(n373), .B1(n372), .B2(n370), .C1(n373), .C2(
        n370), .ZN(p8_C[66]) );
  XNOR2_X1 U419 ( .A(n370), .B(n371), .ZN(p8_S[66]) );
  AOI22_X1 U565 ( .A1(B2[6]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_19_), .ZN(n518) );
  OAI221_X1 U564 ( .B1(B2[5]), .B2(n422), .C1(p8_minus_A_shifted_18_), .C2(
        n423), .A(n518), .ZN(n506) );
  AOI22_X1 U563 ( .A1(B2[4]), .A2(n344), .B1(n345), .B2(p8_minus_A_shifted_17_), .ZN(n517) );
  OAI221_X1 U562 ( .B1(B2[3]), .B2(n341), .C1(p8_minus_A_shifted_16_), .C2(
        n342), .A(n517), .ZN(n507) );
  AOI222_X1 U547 ( .A1(p8_muxs_out_1__15_), .A2(n506), .B1(p8_muxs_out_1__15_), 
        .B2(n507), .C1(n506), .C2(n507), .ZN(n376) );
  XNOR2_X1 U561 ( .A(n506), .B(n507), .ZN(n516) );
  XNOR2_X1 U560 ( .A(p8_muxs_out_1__15_), .B(n516), .ZN(n503) );
  NOR2_X1 U777 ( .A1(reg3_reg[1]), .A2(n2797), .ZN(n560) );
  AOI22_X1 U605 ( .A1(B2[13]), .A2(n560), .B1(reg3_reg[1]), .B2(
        p8_minus_A_shifted_38_), .ZN(n543) );
  NOR2_X1 U588 ( .A1(p8_muxs_out_1__14_), .A2(n543), .ZN(n513) );
  XNOR2_X1 U587 ( .A(p8_muxs_out_1__15_), .B(p8_muxs_out_3__15_), .ZN(n542) );
  XNOR2_X1 U586 ( .A(n542), .B(p8_muxs_out_2__15_), .ZN(n514) );
  AOI22_X1 U602 ( .A1(B2[6]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_19_), .ZN(n559) );
  OAI221_X1 U601 ( .B1(B2[5]), .B2(n437), .C1(p8_minus_A_shifted_18_), .C2(
        n438), .A(n559), .ZN(n544) );
  AOI222_X1 U589 ( .A1(p8_muxs_out_3__14_), .A2(p8_muxs_out_2__14_), .B1(
        p8_muxs_out_3__14_), .B2(n544), .C1(p8_muxs_out_2__14_), .C2(n544), 
        .ZN(n515) );
  AOI222_X1 U559 ( .A1(n513), .A2(n514), .B1(n513), .B2(n515), .C1(n514), .C2(
        n515), .ZN(n504) );
  XNOR2_X1 U553 ( .A(n496), .B(n493), .ZN(n509) );
  XNOR2_X1 U550 ( .A(n509), .B(n494), .ZN(n505) );
  AOI222_X1 U546 ( .A1(n503), .A2(n504), .B1(n503), .B2(n505), .C1(n504), .C2(
        n505), .ZN(n377) );
  XNOR2_X1 U530 ( .A(n492), .B(n491), .ZN(n374) );
  AOI222_X1 U529 ( .A1(n376), .A2(n377), .B1(n376), .B2(n374), .C1(n377), .C2(
        n374), .ZN(p8_C[65]) );
  XNOR2_X1 U421 ( .A(n374), .B(n375), .ZN(p8_S[65]) );
  AOI22_X1 U583 ( .A1(B2[5]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_18_), .ZN(n540) );
  OAI221_X1 U582 ( .B1(B2[4]), .B2(n422), .C1(p8_minus_A_shifted_17_), .C2(
        n423), .A(n540), .ZN(n522) );
  AOI22_X1 U581 ( .A1(B2[3]), .A2(n344), .B1(n345), .B2(p8_minus_A_shifted_16_), .ZN(n539) );
  OAI221_X1 U580 ( .B1(B2[2]), .B2(n341), .C1(p8_minus_A_shifted_15_), .C2(
        n342), .A(n539), .ZN(n523) );
  AOI22_X1 U578 ( .A1(B2[7]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_20_), .ZN(n538) );
  OAI221_X1 U577 ( .B1(B2[6]), .B2(n437), .C1(p8_minus_A_shifted_19_), .C2(
        n438), .A(n538), .ZN(n524) );
  AOI222_X1 U567 ( .A1(n522), .A2(n523), .B1(n522), .B2(n524), .C1(n523), .C2(
        n524), .ZN(n380) );
  XNOR2_X1 U579 ( .A(n522), .B(n523), .ZN(n537) );
  XNOR2_X1 U576 ( .A(n537), .B(n524), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n515), .B(n541), .ZN(n520) );
  NAND2_X1 U773 ( .A1(reg3_reg[1]), .A2(n2797), .ZN(n576) );
  NAND2_X1 U775 ( .A1(reg3_reg[0]), .A2(reg3_reg[1]), .ZN(n594) );
  AOI22_X1 U627 ( .A1(B2[13]), .A2(n560), .B1(n578), .B2(
        p8_minus_A_shifted_38_), .ZN(n577) );
  OAI21_X1 U626 ( .B1(B2[12]), .B2(n576), .A(n577), .ZN(n575) );
  NAND2_X1 U625 ( .A1(n575), .A2(p8_muxs_out_1__13_), .ZN(n534) );
  XNOR2_X1 U603 ( .A(p8_muxs_out_3__14_), .B(p8_muxs_out_2__14_), .ZN(n558) );
  OAI222_X1 U574 ( .A1(n534), .A2(n535), .B1(n534), .B2(n536), .C1(n535), .C2(
        n536), .ZN(n521) );
  AOI222_X1 U566 ( .A1(n519), .A2(n520), .B1(n519), .B2(n521), .C1(n520), .C2(
        n521), .ZN(n379) );
  XNOR2_X1 U558 ( .A(n503), .B(n504), .ZN(n508) );
  AOI222_X1 U548 ( .A1(n380), .A2(n379), .B1(n380), .B2(n381), .C1(n379), .C2(
        n381), .ZN(p8_C[64]) );
  XNOR2_X1 U423 ( .A(n378), .B(n379), .ZN(p8_S[64]) );
  XNOR2_X1 U575 ( .A(n520), .B(n519), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n535), .B(n536), .ZN(n557) );
  AOI22_X1 U632 ( .A1(B2[5]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_18_), .ZN(n580) );
  OAI221_X1 U631 ( .B1(B2[4]), .B2(n437), .C1(p8_minus_A_shifted_17_), .C2(
        n438), .A(n580), .ZN(n564) );
  AOI222_X1 U612 ( .A1(p8_muxs_out_2__13_), .A2(p8_muxs_out_3__13_), .B1(
        p8_muxs_out_2__13_), .B2(n564), .C1(p8_muxs_out_3__13_), .C2(n564), 
        .ZN(n527) );
  AOI22_X1 U611 ( .A1(B2[1]), .A2(n342), .B1(n341), .B2(p8_minus_A_shifted_14_), .ZN(n563) );
  AOI221_X1 U610 ( .B1(n344), .B2(B2[2]), .C1(n345), .C2(
        p8_minus_A_shifted_15_), .A(n563), .ZN(n528) );
  XNOR2_X1 U609 ( .A(n527), .B(n528), .ZN(n561) );
  AOI22_X1 U608 ( .A1(B2[4]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_17_), .ZN(n562) );
  OAI221_X1 U607 ( .B1(B2[3]), .B2(n422), .C1(p8_minus_A_shifted_16_), .C2(
        n423), .A(n562), .ZN(n529) );
  XNOR2_X1 U606 ( .A(n561), .B(n529), .ZN(n531) );
  XNOR2_X1 U629 ( .A(p8_muxs_out_2__13_), .B(n579), .ZN(n554) );
  OAI21_X1 U624 ( .B1(n575), .B2(p8_muxs_out_1__13_), .A(n534), .ZN(n555) );
  OAI222_X1 U654 ( .A1(B2[12]), .A2(n594), .B1(p8_minus_A_shifted_25_), .B2(
        n595), .C1(B2[11]), .C2(n576), .ZN(n593) );
  NAND2_X1 U653 ( .A1(n593), .A2(p8_muxs_out_1__12_), .ZN(n556) );
  AOI222_X1 U596 ( .A1(n554), .A2(n555), .B1(n554), .B2(n556), .C1(n555), .C2(
        n556), .ZN(n532) );
  AOI222_X1 U572 ( .A1(n530), .A2(n531), .B1(n530), .B2(n532), .C1(n531), .C2(
        n532), .ZN(n385) );
  OAI222_X1 U570 ( .A1(n526), .A2(n527), .B1(n526), .B2(n528), .C1(n527), .C2(
        n528), .ZN(n525) );
  AOI222_X1 U568 ( .A1(n384), .A2(n385), .B1(n384), .B2(n382), .C1(n385), .C2(
        n382), .ZN(p8_C[63]) );
  XNOR2_X1 U425 ( .A(n382), .B(n383), .ZN(p8_S[63]) );
  XNOR2_X1 U595 ( .A(n553), .B(n532), .ZN(n388) );
  XNOR2_X1 U623 ( .A(n554), .B(n555), .ZN(n574) );
  AOI22_X1 U659 ( .A1(B2[4]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_17_), .ZN(n597) );
  OAI221_X1 U658 ( .B1(B2[3]), .B2(n437), .C1(p8_minus_A_shifted_16_), .C2(
        n438), .A(n597), .ZN(n587) );
  AOI222_X1 U645 ( .A1(p8_muxs_out_2__12_), .A2(p8_muxs_out_3__12_), .B1(
        p8_muxs_out_2__12_), .B2(n587), .C1(p8_muxs_out_3__12_), .C2(n587), 
        .ZN(n547) );
  AOI22_X1 U639 ( .A1(B2[0]), .A2(n342), .B1(n341), .B2(p8_minus_A_shifted_13_), .ZN(n583) );
  AOI221_X1 U638 ( .B1(n344), .B2(B2[1]), .C1(n345), .C2(
        p8_minus_A_shifted_14_), .A(n583), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n547), .B(n548), .ZN(n581) );
  AOI22_X1 U636 ( .A1(B2[3]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_16_), .ZN(n582) );
  OAI221_X1 U635 ( .B1(B2[2]), .B2(n422), .C1(p8_minus_A_shifted_15_), .C2(
        n423), .A(n582), .ZN(n549) );
  XNOR2_X1 U634 ( .A(n581), .B(n549), .ZN(n551) );
  XNOR2_X1 U656 ( .A(p8_muxs_out_2__12_), .B(n596), .ZN(n571) );
  OAI21_X1 U652 ( .B1(n593), .B2(p8_muxs_out_1__12_), .A(n556), .ZN(n572) );
  AOI22_X1 U678 ( .A1(n617), .A2(p8_minus_A_shifted_23_), .B1(n560), .B2(
        B2[11]), .ZN(n616) );
  OAI21_X1 U677 ( .B1(B2[11]), .B2(n594), .A(n616), .ZN(n615) );
  NAND2_X1 U676 ( .A1(p8_muxs_out_1__11_), .A2(n615), .ZN(n573) );
  AOI222_X1 U620 ( .A1(n571), .A2(n572), .B1(n571), .B2(n573), .C1(n572), .C2(
        n573), .ZN(n552) );
  AOI222_X1 U594 ( .A1(n550), .A2(n551), .B1(n550), .B2(n552), .C1(n551), .C2(
        n552), .ZN(n389) );
  OAI222_X1 U592 ( .A1(n546), .A2(n547), .B1(n546), .B2(n548), .C1(n547), .C2(
        n548), .ZN(n545) );
  AOI222_X1 U590 ( .A1(n388), .A2(n389), .B1(n388), .B2(n386), .C1(n389), .C2(
        n386), .ZN(p8_C[62]) );
  XNOR2_X1 U427 ( .A(n386), .B(n387), .ZN(p8_S[62]) );
  XNOR2_X1 U619 ( .A(n570), .B(n552), .ZN(n392) );
  AOI22_X1 U665 ( .A1(B2[2]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_15_), .ZN(n601) );
  OAI221_X1 U664 ( .B1(B2[1]), .B2(n422), .C1(p8_minus_A_shifted_14_), .C2(
        n423), .A(n601), .ZN(n565) );
  NOR2_X1 U662 ( .A1(n584), .A2(p8_minus_A_shifted_13_), .ZN(n598) );
  XNOR2_X1 U651 ( .A(n571), .B(n572), .ZN(n592) );
  OAI21_X1 U675 ( .B1(p8_muxs_out_1__11_), .B2(n615), .A(n573), .ZN(n602) );
  AOI22_X1 U702 ( .A1(n617), .A2(p8_minus_A_shifted_22_), .B1(n560), .B2(
        B2[10]), .ZN(n630) );
  OAI21_X1 U701 ( .B1(B2[10]), .B2(n594), .A(n630), .ZN(n629) );
  NAND2_X1 U700 ( .A1(p8_muxs_out_1__10_), .A2(n629), .ZN(n604) );
  AOI222_X1 U666 ( .A1(n602), .A2(n603), .B1(n602), .B2(n604), .C1(n603), .C2(
        n604), .ZN(n569) );
  AOI222_X1 U618 ( .A1(n567), .A2(n568), .B1(n567), .B2(n569), .C1(n568), .C2(
        n569), .ZN(n393) );
  OAI221_X1 U615 ( .B1(B2[0]), .B2(n430), .C1(p8_minus_A_shifted_13_), .C2(
        n429), .A(n341), .ZN(n566) );
  AOI222_X1 U614 ( .A1(n565), .A2(reg3_reg[13]), .B1(n565), .B2(n566), .C1(
        reg3_reg[13]), .C2(n566), .ZN(n390) );
  AOI222_X1 U613 ( .A1(n392), .A2(n393), .B1(n392), .B2(n390), .C1(n393), .C2(
        n390), .ZN(p8_C[61]) );
  XNOR2_X1 U429 ( .A(n390), .B(n391), .ZN(p8_S[61]) );
  AOI22_X1 U689 ( .A1(B2[1]), .A2(n425), .B1(n426), .B2(p8_minus_A_shifted_14_), .ZN(n621) );
  OAI221_X1 U688 ( .B1(B2[0]), .B2(n422), .C1(p8_minus_A_shifted_13_), .C2(
        n423), .A(n621), .ZN(n605) );
  AOI22_X1 U685 ( .A1(B2[3]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_16_), .ZN(n620) );
  OAI221_X1 U684 ( .B1(B2[2]), .B2(n437), .C1(p8_minus_A_shifted_15_), .C2(
        n438), .A(n620), .ZN(n606) );
  AOI222_X1 U667 ( .A1(n605), .A2(p8_muxs_out_3__11_), .B1(n605), .B2(n606), 
        .C1(p8_muxs_out_3__11_), .C2(n606), .ZN(n396) );
  XNOR2_X1 U648 ( .A(n569), .B(n591), .ZN(n397) );
  XNOR2_X1 U687 ( .A(n605), .B(p8_muxs_out_3__11_), .ZN(n619) );
  XNOR2_X1 U683 ( .A(n619), .B(n606), .ZN(n588) );
  AOI22_X1 U680 ( .A1(p8_muxs_out_2__11_), .A2(n618), .B1(n604), .B2(n603), 
        .ZN(n614) );
  XNOR2_X1 U674 ( .A(n614), .B(n602), .ZN(n589) );
  OAI21_X1 U699 ( .B1(p8_muxs_out_1__10_), .B2(n629), .A(n604), .ZN(n625) );
  AOI222_X1 U693 ( .A1(n623), .A2(n624), .B1(n623), .B2(n625), .C1(n624), .C2(
        n625), .ZN(n590) );
  AOI222_X1 U647 ( .A1(n588), .A2(n589), .B1(n588), .B2(n590), .C1(n589), .C2(
        n590), .ZN(n394) );
  AOI222_X1 U646 ( .A1(n396), .A2(n397), .B1(n396), .B2(n394), .C1(n397), .C2(
        n394), .ZN(p8_C[60]) );
  AOI22_X1 U711 ( .A1(B2[2]), .A2(n446), .B1(n447), .B2(p8_minus_A_shifted_15_), .ZN(n631) );
  OAI221_X1 U710 ( .B1(B2[1]), .B2(n437), .C1(p8_minus_A_shifted_14_), .C2(
        n438), .A(n631), .ZN(n608) );
  NOR2_X1 U707 ( .A1(n622), .A2(p8_minus_A_shifted_13_), .ZN(n609) );
  XNOR2_X1 U672 ( .A(n590), .B(n613), .ZN(n400) );
  AOI22_X1 U703 ( .A1(p8_muxs_out_2__10_), .A2(p8_muxs_out_3__10_), .B1(n624), 
        .B2(n623), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(n625), .ZN(n611) );
  NOR2_X1 U727 ( .A1(B2[8]), .A2(n576), .ZN(n646) );
  AOI221_X1 U726 ( .B1(B2[9]), .B2(n560), .C1(p8_minus_A_shifted_22_), .C2(
        n578), .A(n646), .ZN(n634) );
  AOI222_X1 U713 ( .A1(n632), .A2(n633), .B1(n632), .B2(n634), .C1(n633), .C2(
        n634), .ZN(n612) );
  AOI222_X1 U671 ( .A1(n610), .A2(n611), .B1(n610), .B2(n612), .C1(n611), .C2(
        n612), .ZN(n401) );
  AOI22_X1 U729 ( .A1(p8_muxs_out_1__9_), .A2(p8_muxs_out_2__9_), .B1(n633), 
        .B2(n632), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(n634), .ZN(n635) );
  AOI22_X1 U723 ( .A1(B2[0]), .A2(n438), .B1(n437), .B2(p8_minus_A_shifted_13_), .ZN(n644) );
  OAI221_X1 U721 ( .B1(n641), .B2(p8_minus_A_shifted_14_), .C1(n642), .C2(
        B2[1]), .A(n643), .ZN(n626) );
  AOI22_X1 U750 ( .A1(B2[8]), .A2(n560), .B1(n578), .B2(p8_minus_A_shifted_21_), .ZN(n656) );
  OAI21_X1 U749 ( .B1(B2[7]), .B2(n576), .A(n656), .ZN(n640) );
  AOI222_X1 U718 ( .A1(p8_muxs_out_1__8_), .A2(p8_muxs_out_2__8_), .B1(
        p8_muxs_out_1__8_), .B2(n640), .C1(p8_muxs_out_2__8_), .C2(n640), .ZN(
        n638) );
  AOI222_X1 U714 ( .A1(n635), .A2(n636), .B1(n635), .B2(n637), .C1(n636), .C2(
        n637), .ZN(n404) );
  XNOR2_X1 U696 ( .A(n612), .B(n627), .ZN(n405) );
  NAND2_X1 U695 ( .A1(p8_muxs_out_3__9_), .A2(n626), .ZN(n402) );
  XNOR2_X1 U719 ( .A(n635), .B(n636), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(n638), .ZN(n406) );
  OAI221_X1 U739 ( .B1(n641), .B2(p8_minus_A_shifted_13_), .C1(n642), .C2(
        B2[0]), .A(n437), .ZN(n647) );
  AOI22_X1 U763 ( .A1(B2[7]), .A2(n595), .B1(n594), .B2(p8_minus_A_shifted_20_), .ZN(n662) );
  AOI21_X1 U762 ( .B1(n617), .B2(p8_minus_A_shifted_19_), .A(n662), .ZN(n660)
         );
  NOR2_X1 U760 ( .A1(n660), .A2(n2856), .ZN(n649) );
  XNOR2_X1 U752 ( .A(p8_muxs_out_2__8_), .B(p8_muxs_out_1__8_), .ZN(n655) );
  XNOR2_X1 U748 ( .A(n655), .B(n640), .ZN(n650) );
  AOI222_X1 U733 ( .A1(n648), .A2(n649), .B1(n648), .B2(n650), .C1(n649), .C2(
        n650), .ZN(n408) );
  NAND2_X1 U732 ( .A1(p8_muxs_out_3__8_), .A2(n647), .ZN(n409) );
  XNOR2_X1 U736 ( .A(n650), .B(n653), .ZN(n410) );
  NOR2_X1 U772 ( .A1(B2[5]), .A2(n576), .ZN(n665) );
  AOI221_X1 U771 ( .B1(B2[6]), .B2(n560), .C1(p8_minus_A_shifted_19_), .C2(
        n578), .A(n665), .ZN(n658) );
  NOR2_X1 U757 ( .A1(n658), .A2(n659), .ZN(n651) );
  AOI22_X1 U440 ( .A1(reg3_reg[9]), .A2(n412), .B1(n413), .B2(n2788), .ZN(n411) );
  XNOR2_X1 U439 ( .A(n410), .B(n411), .ZN(p8_S[56]) );
  XNOR2_X1 U770 ( .A(p8_muxs_out_1__6_), .B(n658), .ZN(n664) );
  NAND2_X1 U769 ( .A1(n664), .A2(p8_muxs_out_2__6_), .ZN(n418) );
  AOI222_X1 U753 ( .A1(n416), .A2(n419), .B1(n416), .B2(n418), .C1(n419), .C2(
        n418), .ZN(p8_C[55]) );
  AOI22_X1 U443 ( .A1(p8_muxs_out_3__7_), .A2(n417), .B1(n418), .B2(n419), 
        .ZN(n415) );
  XNOR2_X1 U442 ( .A(n415), .B(n416), .ZN(p8_S[55]) );
  OAI21_X1 U768 ( .B1(n664), .B2(p8_muxs_out_2__6_), .A(n418), .ZN(n420) );
  NOR2_X1 U767 ( .A1(n663), .A2(n420), .ZN(p8_C[54]) );
  XNOR2_X1 U445 ( .A(p8_muxs_out_3__6_), .B(n420), .ZN(p8_S[54]) );
  AOI222_X1 U668 ( .A1(n400), .A2(n401), .B1(n400), .B2(n398), .C1(n401), .C2(
        n398), .ZN(p8_C[59]) );
  XNOR2_X1 U431 ( .A(n394), .B(n395), .ZN(p8_S[60]) );
  OAI21_X1 U267 ( .B1(reg4_reg[11]), .B2(reg4_reg[12]), .A(n15), .ZN(n260) );
  AOI22_X1 U287 ( .A1(reg4_reg[11]), .A2(n2803), .B1(reg4_reg[12]), .B2(n2787), 
        .ZN(n258) );
  AOI22_X1 U23 ( .A1(B3[13]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_38_), 
        .ZN(n16) );
  OAI221_X1 U22 ( .B1(B3[12]), .B2(n14), .C1(p9_minus_A_shifted_25_), .C2(n15), 
        .A(n16), .ZN(p9_final_product2_26_) );
  AOI22_X1 U71 ( .A1(B3[12]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_25_), 
        .ZN(n95) );
  OAI221_X1 U70 ( .B1(B3[11]), .B2(n14), .C1(n3152), .C2(n15), .A(n95), .ZN(
        p9_C[72]) );
  OAI21_X1 U332 ( .B1(reg4_reg[9]), .B2(reg4_reg[10]), .A(n97), .ZN(n296) );
  AOI22_X1 U86 ( .A1(B3[12]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_25_), 
        .ZN(n114) );
  OAI221_X1 U85 ( .B1(B3[11]), .B2(n96), .C1(n3152), .C2(n97), .A(n114), .ZN(
        n105) );
  OAI21_X1 U370 ( .B1(reg4_reg[8]), .B2(p9_Partial_products_sum_add_23_B_0_), 
        .A(n112), .ZN(n328) );
  AOI22_X1 U96 ( .A1(B3[13]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_38_), .ZN(n113) );
  OAI221_X1 U84 ( .B1(B3[13]), .B2(n111), .C1(p9_minus_A_shifted_38_), .C2(
        n112), .A(n113), .ZN(n108) );
  AOI22_X1 U82 ( .A1(B3[10]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_23_), 
        .ZN(n110) );
  OAI221_X1 U81 ( .B1(B3[9]), .B2(n14), .C1(p9_minus_A_shifted_22_), .C2(n15), 
        .A(n110), .ZN(n107) );
  AOI222_X1 U77 ( .A1(n105), .A2(n106), .B1(n105), .B2(n107), .C1(n106), .C2(
        n107), .ZN(n23) );
  AOI22_X1 U76 ( .A1(B3[11]), .A2(n103), .B1(n104), .B2(n3152), .ZN(n102) );
  AOI221_X1 U75 ( .B1(B3[10]), .B2(n20), .C1(p9_minus_A_shifted_23_), .C2(n101), .A(n102), .ZN(n24) );
  AOI22_X1 U74 ( .A1(B3[13]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_38_), 
        .ZN(n98) );
  OAI221_X1 U73 ( .B1(B3[12]), .B2(n96), .C1(p9_minus_A_shifted_25_), .C2(n97), 
        .A(n98), .ZN(n21) );
  AOI222_X1 U72 ( .A1(n23), .A2(n24), .B1(n23), .B2(n21), .C1(n24), .C2(n21), 
        .ZN(p9_C[71]) );
  XNOR2_X1 U26 ( .A(n21), .B(n22), .ZN(p9_S[71]) );
  OAI221_X1 U95 ( .B1(B3[12]), .B2(n111), .C1(p9_minus_A_shifted_25_), .C2(
        n112), .A(n113), .ZN(n27) );
  AOI22_X1 U94 ( .A1(B3[11]), .A2(n99), .B1(n100), .B2(n3152), .ZN(n119) );
  OAI221_X1 U93 ( .B1(B3[10]), .B2(n96), .C1(p9_minus_A_shifted_23_), .C2(n97), 
        .A(n119), .ZN(n115) );
  AOI22_X1 U117 ( .A1(B3[12]), .A2(n120), .B1(n121), .B2(
        p9_minus_A_shifted_25_), .ZN(n139) );
  OAI221_X1 U116 ( .B1(B3[11]), .B2(n111), .C1(n3152), .C2(n112), .A(n139), 
        .ZN(n122) );
  AOI22_X1 U114 ( .A1(B3[10]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_23_), .ZN(n138) );
  OAI221_X1 U113 ( .B1(B3[9]), .B2(n96), .C1(p9_minus_A_shifted_22_), .C2(n97), 
        .A(n138), .ZN(n123) );
  AOI222_X1 U97 ( .A1(n122), .A2(n123), .B1(n122), .B2(n124), .C1(n123), .C2(
        n124), .ZN(n117) );
  AOI222_X1 U87 ( .A1(n115), .A2(n30), .B1(n115), .B2(n116), .C1(n30), .C2(
        n116), .ZN(n26) );
  XNOR2_X1 U83 ( .A(n105), .B(n108), .ZN(n109) );
  XNOR2_X1 U80 ( .A(n109), .B(n107), .ZN(n29) );
  AOI222_X1 U79 ( .A1(n30), .A2(n26), .B1(n30), .B2(n29), .C1(n26), .C2(n29), 
        .ZN(p9_C[70]) );
  AOI22_X1 U29 ( .A1(n27), .A2(n28), .B1(n29), .B2(n30), .ZN(n25) );
  XNOR2_X1 U28 ( .A(n25), .B(n26), .ZN(p9_S[70]) );
  XNOR2_X1 U115 ( .A(p9_muxs_out_3__20_), .B(n122), .ZN(n137) );
  AOI22_X1 U111 ( .A1(B3[8]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_21_), 
        .ZN(n136) );
  OAI221_X1 U110 ( .B1(B3[7]), .B2(n14), .C1(p9_minus_A_shifted_20_), .C2(n15), 
        .A(n136), .ZN(n127) );
  AOI22_X1 U127 ( .A1(B3[8]), .A2(n97), .B1(n96), .B2(p9_minus_A_shifted_21_), 
        .ZN(n146) );
  AOI221_X1 U126 ( .B1(n99), .B2(B3[9]), .C1(n100), .C2(p9_minus_A_shifted_22_), .A(n146), .ZN(n133) );
  AOI22_X1 U130 ( .A1(B3[11]), .A2(n120), .B1(n121), .B2(n3152), .ZN(n147) );
  OAI221_X1 U129 ( .B1(B3[10]), .B2(n111), .C1(p9_minus_A_shifted_23_), .C2(
        n112), .A(n147), .ZN(n135) );
  AOI222_X1 U107 ( .A1(p9_muxs_out_3__19_), .A2(n133), .B1(p9_muxs_out_3__19_), 
        .B2(n134), .C1(n133), .C2(n134), .ZN(n128) );
  AOI222_X1 U101 ( .A1(n126), .A2(n127), .B1(n126), .B2(n128), .C1(n127), .C2(
        n128), .ZN(n33) );
  AOI22_X1 U100 ( .A1(B3[9]), .A2(n103), .B1(n104), .B2(p9_minus_A_shifted_22_), .ZN(n125) );
  AOI221_X1 U99 ( .B1(B3[8]), .B2(n20), .C1(p9_minus_A_shifted_21_), .C2(n101), 
        .A(n125), .ZN(n34) );
  XNOR2_X1 U91 ( .A(n117), .B(n118), .ZN(n31) );
  AOI222_X1 U90 ( .A1(n33), .A2(n34), .B1(n33), .B2(n31), .C1(n34), .C2(n31), 
        .ZN(p9_C[69]) );
  XNOR2_X1 U31 ( .A(n31), .B(n32), .ZN(p9_S[69]) );
  XNOR2_X1 U106 ( .A(n132), .B(n128), .ZN(n35) );
  XNOR2_X1 U128 ( .A(p9_muxs_out_3__19_), .B(n135), .ZN(n145) );
  AOI22_X1 U147 ( .A1(B3[8]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_21_), 
        .ZN(n160) );
  OAI221_X1 U146 ( .B1(B3[7]), .B2(n96), .C1(p9_minus_A_shifted_20_), .C2(n97), 
        .A(n160), .ZN(n150) );
  AOI22_X1 U144 ( .A1(B3[6]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_19_), 
        .ZN(n159) );
  OAI221_X1 U143 ( .B1(B3[5]), .B2(n14), .C1(p9_minus_A_shifted_18_), .C2(n15), 
        .A(n159), .ZN(n151) );
  AOI222_X1 U135 ( .A1(p9_muxs_out_2__17_), .A2(n150), .B1(p9_muxs_out_2__17_), 
        .B2(n151), .C1(n150), .C2(n151), .ZN(n130) );
  AOI22_X1 U151 ( .A1(B3[10]), .A2(n120), .B1(n121), .B2(
        p9_minus_A_shifted_23_), .ZN(n162) );
  OAI221_X1 U150 ( .B1(B3[9]), .B2(n111), .C1(p9_minus_A_shifted_22_), .C2(
        n112), .A(n162), .ZN(n148) );
  AOI222_X1 U133 ( .A1(p9_muxs_out_3__18_), .A2(n148), .B1(p9_muxs_out_3__18_), 
        .B2(n149), .C1(n148), .C2(n149), .ZN(n131) );
  OAI222_X1 U104 ( .A1(n129), .A2(n130), .B1(n129), .B2(n131), .C1(n130), .C2(
        n131), .ZN(n37) );
  AOI222_X1 U102 ( .A1(n35), .A2(n39), .B1(n35), .B2(n38), .C1(n39), .C2(n38), 
        .ZN(p9_C[68]) );
  AOI22_X1 U34 ( .A1(p9_muxs_out_3__19_), .A2(n37), .B1(n38), .B2(n39), .ZN(
        n36) );
  XNOR2_X1 U33 ( .A(n35), .B(n36), .ZN(p9_S[68]) );
  XNOR2_X1 U132 ( .A(n130), .B(n131), .ZN(n144) );
  XNOR2_X1 U124 ( .A(n144), .B(n129), .ZN(n40) );
  XNOR2_X1 U145 ( .A(p9_muxs_out_2__17_), .B(n150), .ZN(n158) );
  XNOR2_X1 U142 ( .A(n158), .B(n151), .ZN(n141) );
  AOI222_X1 U168 ( .A1(p9_muxs_out_2__16_), .A2(p9_muxs_out_3__16_), .B1(
        p9_muxs_out_2__16_), .B2(n176), .C1(p9_muxs_out_3__16_), .C2(n176), 
        .ZN(n157) );
  AOI222_X1 U140 ( .A1(p9_muxs_out_2__17_), .A2(n156), .B1(p9_muxs_out_2__17_), 
        .B2(n157), .C1(n156), .C2(n157), .ZN(n142) );
  XNOR2_X1 U148 ( .A(p9_muxs_out_2__18_), .B(n161), .ZN(n143) );
  AOI222_X1 U123 ( .A1(n141), .A2(n142), .B1(n141), .B2(n143), .C1(n142), .C2(
        n143), .ZN(n43) );
  OAI22_X1 U120 ( .A1(p9_minus_A_shifted_20_), .A2(n103), .B1(n104), .B2(B3[7]), .ZN(n140) );
  AOI221_X1 U119 ( .B1(p9_minus_A_shifted_19_), .B2(n101), .C1(B3[6]), .C2(n20), .A(n140), .ZN(n42) );
  AOI222_X1 U118 ( .A1(n40), .A2(n43), .B1(n40), .B2(n42), .C1(n43), .C2(n42), 
        .ZN(p9_C[67]) );
  XNOR2_X1 U36 ( .A(n42), .B(n43), .ZN(n41) );
  AOI22_X1 U165 ( .A1(B3[7]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_20_), 
        .ZN(n174) );
  OAI221_X1 U164 ( .B1(B3[6]), .B2(n96), .C1(p9_minus_A_shifted_19_), .C2(n97), 
        .A(n174), .ZN(n152) );
  AOI22_X1 U163 ( .A1(B3[5]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_18_), 
        .ZN(n173) );
  OAI221_X1 U162 ( .B1(B3[4]), .B2(n14), .C1(p9_minus_A_shifted_17_), .C2(n15), 
        .A(n173), .ZN(n153) );
  AOI22_X1 U161 ( .A1(B3[9]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_22_), .ZN(n172) );
  OAI221_X1 U160 ( .B1(B3[8]), .B2(n111), .C1(p9_minus_A_shifted_21_), .C2(
        n112), .A(n172), .ZN(n154) );
  XNOR2_X1 U159 ( .A(n153), .B(n154), .ZN(n171) );
  XNOR2_X1 U158 ( .A(n152), .B(n171), .ZN(n163) );
  XNOR2_X1 U179 ( .A(p9_muxs_out_3__16_), .B(p9_muxs_out_2__16_), .ZN(n185) );
  XNOR2_X1 U178 ( .A(n185), .B(p9_muxs_out_1__16_), .ZN(n167) );
  AOI222_X1 U175 ( .A1(p9_muxs_out_3__15_), .A2(p9_muxs_out_2__15_), .B1(
        p9_muxs_out_3__15_), .B2(n184), .C1(p9_muxs_out_2__15_), .C2(n184), 
        .ZN(n168) );
  AOI22_X1 U181 ( .A1(B3[8]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_21_), .ZN(n186) );
  OAI221_X1 U180 ( .B1(B3[7]), .B2(n111), .C1(p9_minus_A_shifted_20_), .C2(
        n112), .A(n186), .ZN(n170) );
  AOI222_X1 U155 ( .A1(n167), .A2(n168), .B1(n167), .B2(n169), .C1(n168), .C2(
        n169), .ZN(n165) );
  AOI222_X1 U152 ( .A1(n163), .A2(n164), .B1(n163), .B2(n165), .C1(n164), .C2(
        n165), .ZN(n46) );
  XNOR2_X1 U138 ( .A(n143), .B(n155), .ZN(n47) );
  AOI222_X1 U137 ( .A1(n152), .A2(n153), .B1(n152), .B2(n154), .C1(n153), .C2(
        n154), .ZN(n44) );
  AOI222_X1 U136 ( .A1(n46), .A2(n47), .B1(n46), .B2(n44), .C1(n47), .C2(n44), 
        .ZN(p9_C[66]) );
  XNOR2_X1 U37 ( .A(n44), .B(n45), .ZN(p9_S[66]) );
  AOI22_X1 U189 ( .A1(B3[6]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_19_), 
        .ZN(n192) );
  OAI221_X1 U188 ( .B1(B3[5]), .B2(n96), .C1(p9_minus_A_shifted_18_), .C2(n97), 
        .A(n192), .ZN(n180) );
  AOI22_X1 U187 ( .A1(B3[4]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_17_), 
        .ZN(n191) );
  OAI221_X1 U186 ( .B1(B3[3]), .B2(n14), .C1(p9_minus_A_shifted_16_), .C2(n15), 
        .A(n191), .ZN(n181) );
  AOI222_X1 U171 ( .A1(p9_muxs_out_1__15_), .A2(n180), .B1(p9_muxs_out_1__15_), 
        .B2(n181), .C1(n180), .C2(n181), .ZN(n50) );
  XNOR2_X1 U185 ( .A(n180), .B(n181), .ZN(n190) );
  XNOR2_X1 U184 ( .A(p9_muxs_out_1__15_), .B(n190), .ZN(n177) );
  NOR2_X1 U401 ( .A1(reg4_reg[1]), .A2(n2798), .ZN(n234) );
  AOI22_X1 U229 ( .A1(B3[13]), .A2(n234), .B1(reg4_reg[1]), .B2(
        p9_minus_A_shifted_38_), .ZN(n217) );
  NOR2_X1 U212 ( .A1(p9_muxs_out_1__14_), .A2(n217), .ZN(n187) );
  XNOR2_X1 U211 ( .A(p9_muxs_out_1__15_), .B(p9_muxs_out_3__15_), .ZN(n216) );
  XNOR2_X1 U210 ( .A(n216), .B(p9_muxs_out_2__15_), .ZN(n188) );
  AOI22_X1 U226 ( .A1(B3[6]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_19_), .ZN(n233) );
  OAI221_X1 U225 ( .B1(B3[5]), .B2(n111), .C1(p9_minus_A_shifted_18_), .C2(
        n112), .A(n233), .ZN(n218) );
  AOI222_X1 U213 ( .A1(p9_muxs_out_3__14_), .A2(p9_muxs_out_2__14_), .B1(
        p9_muxs_out_3__14_), .B2(n218), .C1(p9_muxs_out_2__14_), .C2(n218), 
        .ZN(n189) );
  AOI222_X1 U183 ( .A1(n187), .A2(n188), .B1(n187), .B2(n189), .C1(n188), .C2(
        n189), .ZN(n178) );
  XNOR2_X1 U177 ( .A(n170), .B(n167), .ZN(n183) );
  XNOR2_X1 U174 ( .A(n183), .B(n168), .ZN(n179) );
  AOI222_X1 U170 ( .A1(n177), .A2(n178), .B1(n177), .B2(n179), .C1(n178), .C2(
        n179), .ZN(n51) );
  XNOR2_X1 U154 ( .A(n166), .B(n165), .ZN(n48) );
  AOI222_X1 U153 ( .A1(n50), .A2(n51), .B1(n50), .B2(n48), .C1(n51), .C2(n48), 
        .ZN(p9_C[65]) );
  XNOR2_X1 U39 ( .A(n48), .B(n49), .ZN(p9_S[65]) );
  AOI22_X1 U207 ( .A1(B3[5]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_18_), 
        .ZN(n214) );
  OAI221_X1 U206 ( .B1(B3[4]), .B2(n96), .C1(p9_minus_A_shifted_17_), .C2(n97), 
        .A(n214), .ZN(n196) );
  AOI22_X1 U205 ( .A1(B3[3]), .A2(n17), .B1(n18), .B2(p9_minus_A_shifted_16_), 
        .ZN(n213) );
  OAI221_X1 U204 ( .B1(B3[2]), .B2(n14), .C1(p9_minus_A_shifted_15_), .C2(n15), 
        .A(n213), .ZN(n197) );
  AOI22_X1 U202 ( .A1(B3[7]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_20_), .ZN(n212) );
  OAI221_X1 U201 ( .B1(B3[6]), .B2(n111), .C1(p9_minus_A_shifted_19_), .C2(
        n112), .A(n212), .ZN(n198) );
  AOI222_X1 U191 ( .A1(n196), .A2(n197), .B1(n196), .B2(n198), .C1(n197), .C2(
        n198), .ZN(n54) );
  XNOR2_X1 U203 ( .A(n196), .B(n197), .ZN(n211) );
  XNOR2_X1 U200 ( .A(n211), .B(n198), .ZN(n193) );
  XNOR2_X1 U208 ( .A(n189), .B(n215), .ZN(n194) );
  NAND2_X1 U397 ( .A1(reg4_reg[1]), .A2(n2798), .ZN(n250) );
  NAND2_X1 U399 ( .A1(reg4_reg[0]), .A2(reg4_reg[1]), .ZN(n268) );
  AOI22_X1 U251 ( .A1(B3[13]), .A2(n234), .B1(n252), .B2(
        p9_minus_A_shifted_38_), .ZN(n251) );
  OAI21_X1 U250 ( .B1(B3[12]), .B2(n250), .A(n251), .ZN(n249) );
  NAND2_X1 U249 ( .A1(n249), .A2(p9_muxs_out_1__13_), .ZN(n208) );
  XNOR2_X1 U227 ( .A(p9_muxs_out_3__14_), .B(p9_muxs_out_2__14_), .ZN(n232) );
  OAI222_X1 U198 ( .A1(n208), .A2(n209), .B1(n208), .B2(n210), .C1(n209), .C2(
        n210), .ZN(n195) );
  AOI222_X1 U190 ( .A1(n193), .A2(n194), .B1(n193), .B2(n195), .C1(n194), .C2(
        n195), .ZN(n53) );
  XNOR2_X1 U182 ( .A(n177), .B(n178), .ZN(n182) );
  AOI222_X1 U172 ( .A1(n54), .A2(n53), .B1(n54), .B2(n55), .C1(n53), .C2(n55), 
        .ZN(p9_C[64]) );
  XNOR2_X1 U41 ( .A(n52), .B(n53), .ZN(p9_S[64]) );
  XNOR2_X1 U199 ( .A(n194), .B(n193), .ZN(n207) );
  XNOR2_X1 U223 ( .A(n209), .B(n210), .ZN(n231) );
  AOI22_X1 U256 ( .A1(B3[5]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_18_), .ZN(n254) );
  OAI221_X1 U255 ( .B1(B3[4]), .B2(n111), .C1(p9_minus_A_shifted_17_), .C2(
        n112), .A(n254), .ZN(n238) );
  AOI222_X1 U236 ( .A1(p9_muxs_out_2__13_), .A2(p9_muxs_out_3__13_), .B1(
        p9_muxs_out_2__13_), .B2(n238), .C1(p9_muxs_out_3__13_), .C2(n238), 
        .ZN(n201) );
  AOI22_X1 U235 ( .A1(B3[1]), .A2(n15), .B1(n14), .B2(p9_minus_A_shifted_14_), 
        .ZN(n237) );
  AOI221_X1 U234 ( .B1(n17), .B2(B3[2]), .C1(n18), .C2(p9_minus_A_shifted_15_), 
        .A(n237), .ZN(n202) );
  XNOR2_X1 U233 ( .A(n201), .B(n202), .ZN(n235) );
  AOI22_X1 U232 ( .A1(B3[4]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_17_), 
        .ZN(n236) );
  OAI221_X1 U231 ( .B1(B3[3]), .B2(n96), .C1(p9_minus_A_shifted_16_), .C2(n97), 
        .A(n236), .ZN(n203) );
  XNOR2_X1 U230 ( .A(n235), .B(n203), .ZN(n205) );
  XNOR2_X1 U253 ( .A(p9_muxs_out_2__13_), .B(n253), .ZN(n228) );
  OAI21_X1 U248 ( .B1(n249), .B2(p9_muxs_out_1__13_), .A(n208), .ZN(n229) );
  OAI222_X1 U278 ( .A1(B3[12]), .A2(n268), .B1(p9_minus_A_shifted_25_), .B2(
        n269), .C1(B3[11]), .C2(n250), .ZN(n267) );
  NAND2_X1 U277 ( .A1(n267), .A2(p9_muxs_out_1__12_), .ZN(n230) );
  AOI222_X1 U220 ( .A1(n228), .A2(n229), .B1(n228), .B2(n230), .C1(n229), .C2(
        n230), .ZN(n206) );
  AOI222_X1 U196 ( .A1(n204), .A2(n205), .B1(n204), .B2(n206), .C1(n205), .C2(
        n206), .ZN(n59) );
  OAI222_X1 U194 ( .A1(n200), .A2(n201), .B1(n200), .B2(n202), .C1(n201), .C2(
        n202), .ZN(n199) );
  AOI222_X1 U192 ( .A1(n58), .A2(n59), .B1(n58), .B2(n56), .C1(n59), .C2(n56), 
        .ZN(p9_C[63]) );
  XNOR2_X1 U43 ( .A(n56), .B(n57), .ZN(p9_S[63]) );
  XNOR2_X1 U219 ( .A(n227), .B(n206), .ZN(n62) );
  XNOR2_X1 U247 ( .A(n228), .B(n229), .ZN(n248) );
  AOI22_X1 U283 ( .A1(B3[4]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_17_), .ZN(n271) );
  OAI221_X1 U282 ( .B1(B3[3]), .B2(n111), .C1(p9_minus_A_shifted_16_), .C2(
        n112), .A(n271), .ZN(n261) );
  AOI222_X1 U269 ( .A1(p9_muxs_out_2__12_), .A2(p9_muxs_out_3__12_), .B1(
        p9_muxs_out_2__12_), .B2(n261), .C1(p9_muxs_out_3__12_), .C2(n261), 
        .ZN(n221) );
  AOI22_X1 U263 ( .A1(B3[0]), .A2(n15), .B1(n14), .B2(p9_minus_A_shifted_13_), 
        .ZN(n257) );
  AOI221_X1 U262 ( .B1(n17), .B2(B3[1]), .C1(n18), .C2(p9_minus_A_shifted_14_), 
        .A(n257), .ZN(n222) );
  XNOR2_X1 U261 ( .A(n221), .B(n222), .ZN(n255) );
  AOI22_X1 U260 ( .A1(B3[3]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_16_), 
        .ZN(n256) );
  OAI221_X1 U259 ( .B1(B3[2]), .B2(n96), .C1(p9_minus_A_shifted_15_), .C2(n97), 
        .A(n256), .ZN(n223) );
  XNOR2_X1 U258 ( .A(n255), .B(n223), .ZN(n225) );
  XNOR2_X1 U280 ( .A(p9_muxs_out_2__12_), .B(n270), .ZN(n245) );
  OAI21_X1 U276 ( .B1(n267), .B2(p9_muxs_out_1__12_), .A(n230), .ZN(n246) );
  AOI22_X1 U302 ( .A1(n291), .A2(p9_minus_A_shifted_23_), .B1(n234), .B2(
        B3[11]), .ZN(n290) );
  OAI21_X1 U301 ( .B1(B3[11]), .B2(n268), .A(n290), .ZN(n289) );
  NAND2_X1 U300 ( .A1(p9_muxs_out_1__11_), .A2(n289), .ZN(n247) );
  AOI222_X1 U244 ( .A1(n245), .A2(n246), .B1(n245), .B2(n247), .C1(n246), .C2(
        n247), .ZN(n226) );
  AOI222_X1 U218 ( .A1(n224), .A2(n225), .B1(n224), .B2(n226), .C1(n225), .C2(
        n226), .ZN(n63) );
  OAI222_X1 U216 ( .A1(n220), .A2(n221), .B1(n220), .B2(n222), .C1(n221), .C2(
        n222), .ZN(n219) );
  AOI222_X1 U214 ( .A1(n62), .A2(n63), .B1(n62), .B2(n60), .C1(n63), .C2(n60), 
        .ZN(p9_C[62]) );
  XNOR2_X1 U45 ( .A(n60), .B(n61), .ZN(p9_S[62]) );
  XNOR2_X1 U243 ( .A(n244), .B(n226), .ZN(n66) );
  AOI22_X1 U289 ( .A1(B3[2]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_15_), 
        .ZN(n275) );
  OAI221_X1 U288 ( .B1(B3[1]), .B2(n96), .C1(p9_minus_A_shifted_14_), .C2(n97), 
        .A(n275), .ZN(n239) );
  NOR2_X1 U286 ( .A1(n258), .A2(p9_minus_A_shifted_13_), .ZN(n272) );
  XNOR2_X1 U275 ( .A(n245), .B(n246), .ZN(n266) );
  OAI21_X1 U299 ( .B1(p9_muxs_out_1__11_), .B2(n289), .A(n247), .ZN(n276) );
  AOI22_X1 U326 ( .A1(n291), .A2(p9_minus_A_shifted_22_), .B1(n234), .B2(
        B3[10]), .ZN(n304) );
  OAI21_X1 U325 ( .B1(B3[10]), .B2(n268), .A(n304), .ZN(n303) );
  NAND2_X1 U324 ( .A1(p9_muxs_out_1__10_), .A2(n303), .ZN(n278) );
  AOI222_X1 U290 ( .A1(n276), .A2(n277), .B1(n276), .B2(n278), .C1(n277), .C2(
        n278), .ZN(n243) );
  AOI222_X1 U242 ( .A1(n241), .A2(n242), .B1(n241), .B2(n243), .C1(n242), .C2(
        n243), .ZN(n67) );
  OAI221_X1 U239 ( .B1(B3[0]), .B2(n104), .C1(p9_minus_A_shifted_13_), .C2(
        n103), .A(n14), .ZN(n240) );
  AOI222_X1 U238 ( .A1(n239), .A2(reg4_reg[13]), .B1(n239), .B2(n240), .C1(
        reg4_reg[13]), .C2(n240), .ZN(n64) );
  AOI222_X1 U237 ( .A1(n66), .A2(n67), .B1(n66), .B2(n64), .C1(n67), .C2(n64), 
        .ZN(p9_C[61]) );
  XNOR2_X1 U53 ( .A(n64), .B(n65), .ZN(p9_S[61]) );
  AOI22_X1 U313 ( .A1(B3[1]), .A2(n99), .B1(n100), .B2(p9_minus_A_shifted_14_), 
        .ZN(n295) );
  OAI221_X1 U312 ( .B1(B3[0]), .B2(n96), .C1(p9_minus_A_shifted_13_), .C2(n97), 
        .A(n295), .ZN(n279) );
  AOI22_X1 U309 ( .A1(B3[3]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_16_), .ZN(n294) );
  OAI221_X1 U308 ( .B1(B3[2]), .B2(n111), .C1(p9_minus_A_shifted_15_), .C2(
        n112), .A(n294), .ZN(n280) );
  AOI222_X1 U291 ( .A1(n279), .A2(p9_muxs_out_3__11_), .B1(n279), .B2(n280), 
        .C1(p9_muxs_out_3__11_), .C2(n280), .ZN(n70) );
  XNOR2_X1 U272 ( .A(n243), .B(n265), .ZN(n71) );
  XNOR2_X1 U311 ( .A(n279), .B(p9_muxs_out_3__11_), .ZN(n293) );
  XNOR2_X1 U307 ( .A(n293), .B(n280), .ZN(n262) );
  AOI22_X1 U304 ( .A1(p9_muxs_out_2__11_), .A2(n292), .B1(n278), .B2(n277), 
        .ZN(n288) );
  XNOR2_X1 U298 ( .A(n288), .B(n276), .ZN(n263) );
  OAI21_X1 U323 ( .B1(p9_muxs_out_1__10_), .B2(n303), .A(n278), .ZN(n299) );
  AOI222_X1 U317 ( .A1(n297), .A2(n298), .B1(n297), .B2(n299), .C1(n298), .C2(
        n299), .ZN(n264) );
  AOI222_X1 U271 ( .A1(n262), .A2(n263), .B1(n262), .B2(n264), .C1(n263), .C2(
        n264), .ZN(n68) );
  AOI222_X1 U270 ( .A1(n70), .A2(n71), .B1(n70), .B2(n68), .C1(n71), .C2(n68), 
        .ZN(p9_C[60]) );
  AOI22_X1 U335 ( .A1(B3[2]), .A2(n120), .B1(n121), .B2(p9_minus_A_shifted_15_), .ZN(n305) );
  OAI221_X1 U334 ( .B1(B3[1]), .B2(n111), .C1(p9_minus_A_shifted_14_), .C2(
        n112), .A(n305), .ZN(n282) );
  NOR2_X1 U331 ( .A1(n296), .A2(p9_minus_A_shifted_13_), .ZN(n283) );
  XNOR2_X1 U296 ( .A(n264), .B(n287), .ZN(n74) );
  AOI22_X1 U327 ( .A1(p9_muxs_out_2__10_), .A2(p9_muxs_out_3__10_), .B1(n298), 
        .B2(n297), .ZN(n302) );
  XNOR2_X1 U322 ( .A(n302), .B(n299), .ZN(n285) );
  NOR2_X1 U351 ( .A1(B3[8]), .A2(n250), .ZN(n320) );
  AOI221_X1 U350 ( .B1(B3[9]), .B2(n234), .C1(p9_minus_A_shifted_22_), .C2(
        n252), .A(n320), .ZN(n308) );
  AOI222_X1 U337 ( .A1(n306), .A2(n307), .B1(n306), .B2(n308), .C1(n307), .C2(
        n308), .ZN(n286) );
  AOI222_X1 U295 ( .A1(n284), .A2(n285), .B1(n284), .B2(n286), .C1(n285), .C2(
        n286), .ZN(n75) );
  AOI22_X1 U353 ( .A1(p9_muxs_out_1__9_), .A2(p9_muxs_out_2__9_), .B1(n307), 
        .B2(n306), .ZN(n319) );
  XNOR2_X1 U349 ( .A(n319), .B(n308), .ZN(n309) );
  AOI22_X1 U347 ( .A1(B3[0]), .A2(n112), .B1(n111), .B2(p9_minus_A_shifted_13_), .ZN(n318) );
  OAI221_X1 U345 ( .B1(n315), .B2(p9_minus_A_shifted_14_), .C1(n316), .C2(
        B3[1]), .A(n317), .ZN(n300) );
  AOI22_X1 U374 ( .A1(B3[8]), .A2(n234), .B1(n252), .B2(p9_minus_A_shifted_21_), .ZN(n330) );
  OAI21_X1 U373 ( .B1(B3[7]), .B2(n250), .A(n330), .ZN(n314) );
  AOI222_X1 U342 ( .A1(p9_muxs_out_1__8_), .A2(p9_muxs_out_2__8_), .B1(
        p9_muxs_out_1__8_), .B2(n314), .C1(p9_muxs_out_2__8_), .C2(n314), .ZN(
        n312) );
  AOI222_X1 U338 ( .A1(n309), .A2(n310), .B1(n309), .B2(n311), .C1(n310), .C2(
        n311), .ZN(n78) );
  XNOR2_X1 U320 ( .A(n286), .B(n301), .ZN(n79) );
  NAND2_X1 U319 ( .A1(p9_muxs_out_3__9_), .A2(n300), .ZN(n76) );
  XNOR2_X1 U343 ( .A(n309), .B(n310), .ZN(n313) );
  XNOR2_X1 U341 ( .A(n313), .B(n312), .ZN(n80) );
  OAI221_X1 U363 ( .B1(n315), .B2(p9_minus_A_shifted_13_), .C1(n316), .C2(
        B3[0]), .A(n111), .ZN(n321) );
  AOI22_X1 U387 ( .A1(B3[7]), .A2(n269), .B1(n268), .B2(p9_minus_A_shifted_20_), .ZN(n336) );
  AOI21_X1 U386 ( .B1(n291), .B2(p9_minus_A_shifted_19_), .A(n336), .ZN(n334)
         );
  NOR2_X1 U384 ( .A1(n334), .A2(n2857), .ZN(n323) );
  XNOR2_X1 U376 ( .A(p9_muxs_out_2__8_), .B(p9_muxs_out_1__8_), .ZN(n329) );
  XNOR2_X1 U372 ( .A(n329), .B(n314), .ZN(n324) );
  AOI222_X1 U357 ( .A1(n322), .A2(n323), .B1(n322), .B2(n324), .C1(n323), .C2(
        n324), .ZN(n82) );
  NAND2_X1 U356 ( .A1(p9_muxs_out_3__8_), .A2(n321), .ZN(n83) );
  XNOR2_X1 U360 ( .A(n324), .B(n327), .ZN(n84) );
  NOR2_X1 U396 ( .A1(B3[5]), .A2(n250), .ZN(n339) );
  AOI221_X1 U395 ( .B1(B3[6]), .B2(n234), .C1(p9_minus_A_shifted_19_), .C2(
        n252), .A(n339), .ZN(n332) );
  NOR2_X1 U381 ( .A1(n332), .A2(n333), .ZN(n325) );
  AOI22_X1 U64 ( .A1(reg4_reg[9]), .A2(n86), .B1(n87), .B2(n2789), .ZN(n85) );
  XNOR2_X1 U63 ( .A(n84), .B(n85), .ZN(p9_S[56]) );
  XNOR2_X1 U394 ( .A(p9_muxs_out_1__6_), .B(n332), .ZN(n338) );
  NAND2_X1 U393 ( .A1(n338), .A2(p9_muxs_out_2__6_), .ZN(n92) );
  AOI222_X1 U377 ( .A1(n90), .A2(n93), .B1(n90), .B2(n92), .C1(n93), .C2(n92), 
        .ZN(p9_C[55]) );
  AOI22_X1 U67 ( .A1(p9_muxs_out_3__7_), .A2(n91), .B1(n92), .B2(n93), .ZN(n89) );
  XNOR2_X1 U66 ( .A(n89), .B(n90), .ZN(p9_S[55]) );
  OAI21_X1 U392 ( .B1(n338), .B2(p9_muxs_out_2__6_), .A(n92), .ZN(n94) );
  NOR2_X1 U391 ( .A1(n337), .A2(n94), .ZN(p9_C[54]) );
  XNOR2_X1 U69 ( .A(p9_muxs_out_3__6_), .B(n94), .ZN(p9_S[54]) );
  AOI222_X1 U292 ( .A1(n74), .A2(n75), .B1(n74), .B2(n72), .C1(n75), .C2(n72), 
        .ZN(p9_C[59]) );
  XNOR2_X1 U55 ( .A(n68), .B(n69), .ZN(p9_S[60]) );
  OAI21_X1 U1019 ( .B1(reg2_reg[11]), .B2(reg2_reg[12]), .A(n668), .ZN(n912)
         );
  AOI22_X1 U1039 ( .A1(reg2_reg[11]), .A2(n2849), .B1(reg2_reg[12]), .B2(n2791), .ZN(n910) );
  AOI22_X1 U781 ( .A1(B1[13]), .A2(n670), .B1(n671), .B2(
        p7_minus_A_shifted_38_), .ZN(n669) );
  OAI221_X1 U780 ( .B1(B1[12]), .B2(n667), .C1(p7_minus_A_shifted_25_), .C2(
        n668), .A(n669), .ZN(p7_final_product2_26_) );
  AOI22_X1 U823 ( .A1(B1[12]), .A2(n670), .B1(n671), .B2(
        p7_minus_A_shifted_25_), .ZN(n747) );
  OAI221_X1 U822 ( .B1(B1[11]), .B2(n667), .C1(n2984), .C2(n668), .A(n747), 
        .ZN(p7_C[72]) );
  OAI21_X1 U1084 ( .B1(reg2_reg[9]), .B2(reg2_reg[10]), .A(n749), .ZN(n948) );
  AOI22_X1 U838 ( .A1(B1[12]), .A2(n751), .B1(n752), .B2(
        p7_minus_A_shifted_25_), .ZN(n766) );
  OAI221_X1 U837 ( .B1(B1[11]), .B2(n748), .C1(n2984), .C2(n749), .A(n766), 
        .ZN(n757) );
  OAI21_X1 U1122 ( .B1(reg2_reg[8]), .B2(p7_Partial_products_sum_add_23_B_0_), 
        .A(n764), .ZN(n980) );
  AOI22_X1 U848 ( .A1(B1[13]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_38_), .ZN(n765) );
  OAI221_X1 U836 ( .B1(B1[13]), .B2(n763), .C1(p7_minus_A_shifted_38_), .C2(
        n764), .A(n765), .ZN(n760) );
  AOI22_X1 U834 ( .A1(B1[10]), .A2(n670), .B1(n671), .B2(
        p7_minus_A_shifted_23_), .ZN(n762) );
  OAI221_X1 U833 ( .B1(B1[9]), .B2(n667), .C1(p7_minus_A_shifted_22_), .C2(
        n668), .A(n762), .ZN(n759) );
  AOI222_X1 U829 ( .A1(n757), .A2(n758), .B1(n757), .B2(n759), .C1(n758), .C2(
        n759), .ZN(n675) );
  AOI22_X1 U828 ( .A1(B1[11]), .A2(n755), .B1(n756), .B2(n2984), .ZN(n754) );
  AOI221_X1 U827 ( .B1(B1[10]), .B2(n672), .C1(p7_minus_A_shifted_23_), .C2(
        n753), .A(n754), .ZN(n676) );
  AOI22_X1 U826 ( .A1(B1[13]), .A2(n751), .B1(n752), .B2(
        p7_minus_A_shifted_38_), .ZN(n750) );
  OAI221_X1 U825 ( .B1(B1[12]), .B2(n748), .C1(p7_minus_A_shifted_25_), .C2(
        n749), .A(n750), .ZN(n673) );
  AOI222_X1 U824 ( .A1(n675), .A2(n676), .B1(n675), .B2(n673), .C1(n676), .C2(
        n673), .ZN(p7_C[71]) );
  XNOR2_X1 U784 ( .A(n673), .B(n674), .ZN(p7_S[71]) );
  OAI221_X1 U847 ( .B1(B1[12]), .B2(n763), .C1(p7_minus_A_shifted_25_), .C2(
        n764), .A(n765), .ZN(n679) );
  AOI22_X1 U846 ( .A1(B1[11]), .A2(n751), .B1(n752), .B2(n2984), .ZN(n771) );
  OAI221_X1 U845 ( .B1(B1[10]), .B2(n748), .C1(p7_minus_A_shifted_23_), .C2(
        n749), .A(n771), .ZN(n767) );
  AOI22_X1 U869 ( .A1(B1[12]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_25_), .ZN(n791) );
  OAI221_X1 U868 ( .B1(B1[11]), .B2(n763), .C1(n2984), .C2(n764), .A(n791), 
        .ZN(n774) );
  AOI22_X1 U866 ( .A1(B1[10]), .A2(n751), .B1(n752), .B2(
        p7_minus_A_shifted_23_), .ZN(n790) );
  OAI221_X1 U865 ( .B1(B1[9]), .B2(n748), .C1(p7_minus_A_shifted_22_), .C2(
        n749), .A(n790), .ZN(n775) );
  AOI222_X1 U849 ( .A1(n774), .A2(n775), .B1(n774), .B2(n776), .C1(n775), .C2(
        n776), .ZN(n769) );
  AOI222_X1 U839 ( .A1(n767), .A2(n682), .B1(n767), .B2(n768), .C1(n682), .C2(
        n768), .ZN(n678) );
  XNOR2_X1 U835 ( .A(n757), .B(n760), .ZN(n761) );
  XNOR2_X1 U832 ( .A(n761), .B(n759), .ZN(n681) );
  AOI222_X1 U831 ( .A1(n682), .A2(n678), .B1(n682), .B2(n681), .C1(n678), .C2(
        n681), .ZN(p7_C[70]) );
  AOI22_X1 U787 ( .A1(n679), .A2(n680), .B1(n681), .B2(n682), .ZN(n677) );
  XNOR2_X1 U786 ( .A(n677), .B(n678), .ZN(p7_S[70]) );
  XNOR2_X1 U867 ( .A(p7_muxs_out_3__20_), .B(n774), .ZN(n789) );
  AOI22_X1 U863 ( .A1(B1[8]), .A2(n670), .B1(n671), .B2(p7_minus_A_shifted_21_), .ZN(n788) );
  OAI221_X1 U862 ( .B1(B1[7]), .B2(n667), .C1(p7_minus_A_shifted_20_), .C2(
        n668), .A(n788), .ZN(n779) );
  AOI22_X1 U879 ( .A1(B1[8]), .A2(n749), .B1(n748), .B2(p7_minus_A_shifted_21_), .ZN(n798) );
  AOI221_X1 U878 ( .B1(n751), .B2(B1[9]), .C1(n752), .C2(
        p7_minus_A_shifted_22_), .A(n798), .ZN(n785) );
  AOI22_X1 U882 ( .A1(B1[11]), .A2(n772), .B1(n773), .B2(n2984), .ZN(n799) );
  OAI221_X1 U881 ( .B1(B1[10]), .B2(n763), .C1(p7_minus_A_shifted_23_), .C2(
        n764), .A(n799), .ZN(n787) );
  AOI222_X1 U859 ( .A1(p7_muxs_out_3__19_), .A2(n785), .B1(p7_muxs_out_3__19_), 
        .B2(n786), .C1(n785), .C2(n786), .ZN(n780) );
  AOI222_X1 U853 ( .A1(n778), .A2(n779), .B1(n778), .B2(n780), .C1(n779), .C2(
        n780), .ZN(n685) );
  AOI22_X1 U852 ( .A1(B1[9]), .A2(n755), .B1(n756), .B2(p7_minus_A_shifted_22_), .ZN(n777) );
  AOI221_X1 U851 ( .B1(B1[8]), .B2(n672), .C1(p7_minus_A_shifted_21_), .C2(
        n753), .A(n777), .ZN(n686) );
  XNOR2_X1 U843 ( .A(n769), .B(n770), .ZN(n683) );
  AOI222_X1 U842 ( .A1(n685), .A2(n686), .B1(n685), .B2(n683), .C1(n686), .C2(
        n683), .ZN(p7_C[69]) );
  XNOR2_X1 U789 ( .A(n683), .B(n684), .ZN(p7_S[69]) );
  XNOR2_X1 U858 ( .A(n784), .B(n780), .ZN(n687) );
  XNOR2_X1 U880 ( .A(p7_muxs_out_3__19_), .B(n787), .ZN(n797) );
  AOI22_X1 U899 ( .A1(B1[8]), .A2(n751), .B1(n752), .B2(p7_minus_A_shifted_21_), .ZN(n812) );
  OAI221_X1 U898 ( .B1(B1[7]), .B2(n748), .C1(p7_minus_A_shifted_20_), .C2(
        n749), .A(n812), .ZN(n802) );
  AOI22_X1 U896 ( .A1(B1[6]), .A2(n670), .B1(n671), .B2(p7_minus_A_shifted_19_), .ZN(n811) );
  OAI221_X1 U895 ( .B1(B1[5]), .B2(n667), .C1(p7_minus_A_shifted_18_), .C2(
        n668), .A(n811), .ZN(n803) );
  AOI222_X1 U887 ( .A1(p7_muxs_out_2__17_), .A2(n802), .B1(p7_muxs_out_2__17_), 
        .B2(n803), .C1(n802), .C2(n803), .ZN(n782) );
  AOI22_X1 U903 ( .A1(B1[10]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_23_), .ZN(n814) );
  OAI221_X1 U902 ( .B1(B1[9]), .B2(n763), .C1(p7_minus_A_shifted_22_), .C2(
        n764), .A(n814), .ZN(n800) );
  AOI222_X1 U885 ( .A1(p7_muxs_out_3__18_), .A2(n800), .B1(p7_muxs_out_3__18_), 
        .B2(n801), .C1(n800), .C2(n801), .ZN(n783) );
  OAI222_X1 U856 ( .A1(n781), .A2(n782), .B1(n781), .B2(n783), .C1(n782), .C2(
        n783), .ZN(n689) );
  AOI222_X1 U854 ( .A1(n687), .A2(n691), .B1(n687), .B2(n690), .C1(n691), .C2(
        n690), .ZN(p7_C[68]) );
  AOI22_X1 U792 ( .A1(p7_muxs_out_3__19_), .A2(n689), .B1(n690), .B2(n691), 
        .ZN(n688) );
  XNOR2_X1 U791 ( .A(n687), .B(n688), .ZN(p7_S[68]) );
  XNOR2_X1 U884 ( .A(n782), .B(n783), .ZN(n796) );
  XNOR2_X1 U876 ( .A(n796), .B(n781), .ZN(n692) );
  XNOR2_X1 U897 ( .A(p7_muxs_out_2__17_), .B(n802), .ZN(n810) );
  XNOR2_X1 U894 ( .A(n810), .B(n803), .ZN(n793) );
  AOI222_X1 U920 ( .A1(p7_muxs_out_2__16_), .A2(p7_muxs_out_3__16_), .B1(
        p7_muxs_out_2__16_), .B2(n828), .C1(p7_muxs_out_3__16_), .C2(n828), 
        .ZN(n809) );
  AOI222_X1 U892 ( .A1(p7_muxs_out_2__17_), .A2(n808), .B1(p7_muxs_out_2__17_), 
        .B2(n809), .C1(n808), .C2(n809), .ZN(n794) );
  XNOR2_X1 U900 ( .A(p7_muxs_out_2__18_), .B(n813), .ZN(n795) );
  AOI222_X1 U875 ( .A1(n793), .A2(n794), .B1(n793), .B2(n795), .C1(n794), .C2(
        n795), .ZN(n695) );
  OAI22_X1 U872 ( .A1(p7_minus_A_shifted_20_), .A2(n755), .B1(n756), .B2(B1[7]), .ZN(n792) );
  AOI221_X1 U871 ( .B1(p7_minus_A_shifted_19_), .B2(n753), .C1(B1[6]), .C2(
        n672), .A(n792), .ZN(n694) );
  AOI222_X1 U870 ( .A1(n692), .A2(n695), .B1(n692), .B2(n694), .C1(n695), .C2(
        n694), .ZN(p7_C[67]) );
  XNOR2_X1 U794 ( .A(n694), .B(n695), .ZN(n693) );
  AOI22_X1 U917 ( .A1(B1[7]), .A2(n751), .B1(n752), .B2(p7_minus_A_shifted_20_), .ZN(n826) );
  OAI221_X1 U916 ( .B1(B1[6]), .B2(n748), .C1(p7_minus_A_shifted_19_), .C2(
        n749), .A(n826), .ZN(n804) );
  AOI22_X1 U915 ( .A1(B1[5]), .A2(n670), .B1(n671), .B2(p7_minus_A_shifted_18_), .ZN(n825) );
  OAI221_X1 U914 ( .B1(B1[4]), .B2(n667), .C1(p7_minus_A_shifted_17_), .C2(
        n668), .A(n825), .ZN(n805) );
  AOI22_X1 U913 ( .A1(B1[9]), .A2(n772), .B1(n773), .B2(p7_minus_A_shifted_22_), .ZN(n824) );
  OAI221_X1 U912 ( .B1(B1[8]), .B2(n763), .C1(p7_minus_A_shifted_21_), .C2(
        n764), .A(n824), .ZN(n806) );
  XNOR2_X1 U911 ( .A(n805), .B(n806), .ZN(n823) );
  XNOR2_X1 U910 ( .A(n804), .B(n823), .ZN(n815) );
  XNOR2_X1 U931 ( .A(p7_muxs_out_3__16_), .B(p7_muxs_out_2__16_), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n837), .B(p7_muxs_out_1__16_), .ZN(n819) );
  AOI222_X1 U927 ( .A1(p7_muxs_out_3__15_), .A2(p7_muxs_out_2__15_), .B1(
        p7_muxs_out_3__15_), .B2(n836), .C1(p7_muxs_out_2__15_), .C2(n836), 
        .ZN(n820) );
  AOI22_X1 U933 ( .A1(B1[8]), .A2(n772), .B1(n773), .B2(p7_minus_A_shifted_21_), .ZN(n838) );
  OAI221_X1 U932 ( .B1(B1[7]), .B2(n763), .C1(p7_minus_A_shifted_20_), .C2(
        n764), .A(n838), .ZN(n822) );
  AOI222_X1 U907 ( .A1(n819), .A2(n820), .B1(n819), .B2(n821), .C1(n820), .C2(
        n821), .ZN(n817) );
  AOI222_X1 U904 ( .A1(n815), .A2(n816), .B1(n815), .B2(n817), .C1(n816), .C2(
        n817), .ZN(n698) );
  XNOR2_X1 U890 ( .A(n795), .B(n807), .ZN(n699) );
  AOI222_X1 U889 ( .A1(n804), .A2(n805), .B1(n804), .B2(n806), .C1(n805), .C2(
        n806), .ZN(n696) );
  AOI222_X1 U888 ( .A1(n698), .A2(n699), .B1(n698), .B2(n696), .C1(n699), .C2(
        n696), .ZN(p7_C[66]) );
  XNOR2_X1 U795 ( .A(n696), .B(n697), .ZN(p7_S[66]) );
  AOI22_X1 U941 ( .A1(B1[6]), .A2(n751), .B1(n752), .B2(p7_minus_A_shifted_19_), .ZN(n844) );
  OAI221_X1 U940 ( .B1(B1[5]), .B2(n748), .C1(p7_minus_A_shifted_18_), .C2(
        n749), .A(n844), .ZN(n832) );
  AOI22_X1 U939 ( .A1(B1[4]), .A2(n670), .B1(n671), .B2(p7_minus_A_shifted_17_), .ZN(n843) );
  OAI221_X1 U938 ( .B1(B1[3]), .B2(n667), .C1(p7_minus_A_shifted_16_), .C2(
        n668), .A(n843), .ZN(n833) );
  AOI222_X1 U923 ( .A1(p7_muxs_out_1__15_), .A2(n832), .B1(p7_muxs_out_1__15_), 
        .B2(n833), .C1(n832), .C2(n833), .ZN(n702) );
  XNOR2_X1 U937 ( .A(n832), .B(n833), .ZN(n842) );
  XNOR2_X1 U936 ( .A(p7_muxs_out_1__15_), .B(n842), .ZN(n829) );
  NOR2_X1 U1153 ( .A1(reg2_reg[1]), .A2(n2837), .ZN(n886) );
  AOI22_X1 U981 ( .A1(B1[13]), .A2(n886), .B1(reg2_reg[1]), .B2(
        p7_minus_A_shifted_38_), .ZN(n869) );
  NOR2_X1 U964 ( .A1(p7_muxs_out_1__14_), .A2(n869), .ZN(n839) );
  XNOR2_X1 U963 ( .A(p7_muxs_out_1__15_), .B(p7_muxs_out_3__15_), .ZN(n868) );
  XNOR2_X1 U962 ( .A(n868), .B(p7_muxs_out_2__15_), .ZN(n840) );
  AOI22_X1 U978 ( .A1(B1[6]), .A2(n772), .B1(n773), .B2(p7_minus_A_shifted_19_), .ZN(n885) );
  OAI221_X1 U977 ( .B1(B1[5]), .B2(n763), .C1(p7_minus_A_shifted_18_), .C2(
        n764), .A(n885), .ZN(n870) );
  AOI222_X1 U965 ( .A1(p7_muxs_out_3__14_), .A2(p7_muxs_out_2__14_), .B1(
        p7_muxs_out_3__14_), .B2(n870), .C1(p7_muxs_out_2__14_), .C2(n870), 
        .ZN(n841) );
  AOI222_X1 U935 ( .A1(n839), .A2(n840), .B1(n839), .B2(n841), .C1(n840), .C2(
        n841), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n822), .B(n819), .ZN(n835) );
  XNOR2_X1 U926 ( .A(n835), .B(n820), .ZN(n831) );
  AOI222_X1 U922 ( .A1(n829), .A2(n830), .B1(n829), .B2(n831), .C1(n830), .C2(
        n831), .ZN(n703) );
  XNOR2_X1 U906 ( .A(n818), .B(n817), .ZN(n700) );
  AOI222_X1 U905 ( .A1(n702), .A2(n703), .B1(n702), .B2(n700), .C1(n703), .C2(
        n700), .ZN(p7_C[65]) );
  XNOR2_X1 U797 ( .A(n700), .B(n701), .ZN(p7_S[65]) );
  AOI22_X1 U959 ( .A1(B1[5]), .A2(n751), .B1(n752), .B2(p7_minus_A_shifted_18_), .ZN(n866) );
  OAI221_X1 U958 ( .B1(B1[4]), .B2(n748), .C1(p7_minus_A_shifted_17_), .C2(
        n749), .A(n866), .ZN(n848) );
  AOI22_X1 U957 ( .A1(B1[3]), .A2(n670), .B1(n671), .B2(p7_minus_A_shifted_16_), .ZN(n865) );
  OAI221_X1 U956 ( .B1(B1[2]), .B2(n667), .C1(p7_minus_A_shifted_15_), .C2(
        n668), .A(n865), .ZN(n849) );
  AOI22_X1 U954 ( .A1(B1[7]), .A2(n772), .B1(n773), .B2(p7_minus_A_shifted_20_), .ZN(n864) );
  OAI221_X1 U953 ( .B1(B1[6]), .B2(n763), .C1(p7_minus_A_shifted_19_), .C2(
        n764), .A(n864), .ZN(n850) );
  AOI222_X1 U943 ( .A1(n848), .A2(n849), .B1(n848), .B2(n850), .C1(n849), .C2(
        n850), .ZN(n706) );
  XNOR2_X1 U955 ( .A(n848), .B(n849), .ZN(n863) );
  XNOR2_X1 U952 ( .A(n863), .B(n850), .ZN(n845) );
  XNOR2_X1 U960 ( .A(n841), .B(n867), .ZN(n846) );
  NAND2_X1 U1149 ( .A1(reg2_reg[1]), .A2(n2837), .ZN(n902) );
  NAND2_X1 U1151 ( .A1(reg2_reg[0]), .A2(reg2_reg[1]), .ZN(n920) );
  AOI22_X1 U1003 ( .A1(B1[13]), .A2(n886), .B1(n904), .B2(
        p7_minus_A_shifted_38_), .ZN(n903) );
  OAI21_X1 U1002 ( .B1(B1[12]), .B2(n902), .A(n903), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n901), .A2(p7_muxs_out_1__13_), .ZN(n860) );
  XNOR2_X1 U979 ( .A(p7_muxs_out_3__14_), .B(p7_muxs_out_2__14_), .ZN(n884) );
  OAI222_X1 U950 ( .A1(n860), .A2(n861), .B1(n860), .B2(n862), .C1(n861), .C2(
        n862), .ZN(n847) );
  AOI222_X1 U942 ( .A1(n845), .A2(n846), .B1(n845), .B2(n847), .C1(n846), .C2(
        n847), .ZN(n705) );
  XNOR2_X1 U934 ( .A(n829), .B(n830), .ZN(n834) );
  AOI222_X1 U924 ( .A1(n706), .A2(n705), .B1(n706), .B2(n707), .C1(n705), .C2(
        n707), .ZN(p7_C[64]) );
  XNOR2_X1 U799 ( .A(n704), .B(n705), .ZN(p7_S[64]) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n859) );
  XNOR2_X1 U975 ( .A(n861), .B(n862), .ZN(n883) );
  AOI22_X1 U1008 ( .A1(B1[5]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_18_), .ZN(n906) );
  OAI221_X1 U1007 ( .B1(B1[4]), .B2(n763), .C1(p7_minus_A_shifted_17_), .C2(
        n764), .A(n906), .ZN(n890) );
  AOI222_X1 U988 ( .A1(p7_muxs_out_2__13_), .A2(p7_muxs_out_3__13_), .B1(
        p7_muxs_out_2__13_), .B2(n890), .C1(p7_muxs_out_3__13_), .C2(n890), 
        .ZN(n853) );
  AOI22_X1 U987 ( .A1(B1[1]), .A2(n668), .B1(n667), .B2(p7_minus_A_shifted_14_), .ZN(n889) );
  AOI221_X1 U986 ( .B1(n670), .B2(B1[2]), .C1(n671), .C2(
        p7_minus_A_shifted_15_), .A(n889), .ZN(n854) );
  XNOR2_X1 U985 ( .A(n853), .B(n854), .ZN(n887) );
  AOI22_X1 U984 ( .A1(B1[4]), .A2(n751), .B1(n752), .B2(p7_minus_A_shifted_17_), .ZN(n888) );
  OAI221_X1 U983 ( .B1(B1[3]), .B2(n748), .C1(p7_minus_A_shifted_16_), .C2(
        n749), .A(n888), .ZN(n855) );
  XNOR2_X1 U982 ( .A(n887), .B(n855), .ZN(n857) );
  XNOR2_X1 U1005 ( .A(p7_muxs_out_2__13_), .B(n905), .ZN(n880) );
  OAI21_X1 U1000 ( .B1(n901), .B2(p7_muxs_out_1__13_), .A(n860), .ZN(n881) );
  OAI222_X1 U1030 ( .A1(B1[12]), .A2(n920), .B1(p7_minus_A_shifted_25_), .B2(
        n921), .C1(B1[11]), .C2(n902), .ZN(n919) );
  NAND2_X1 U1029 ( .A1(n919), .A2(p7_muxs_out_1__12_), .ZN(n882) );
  AOI222_X1 U972 ( .A1(n880), .A2(n881), .B1(n880), .B2(n882), .C1(n881), .C2(
        n882), .ZN(n858) );
  AOI222_X1 U948 ( .A1(n856), .A2(n857), .B1(n856), .B2(n858), .C1(n857), .C2(
        n858), .ZN(n711) );
  OAI222_X1 U946 ( .A1(n852), .A2(n853), .B1(n852), .B2(n854), .C1(n853), .C2(
        n854), .ZN(n851) );
  AOI222_X1 U944 ( .A1(n710), .A2(n711), .B1(n710), .B2(n708), .C1(n711), .C2(
        n708), .ZN(p7_C[63]) );
  XNOR2_X1 U801 ( .A(n708), .B(n709), .ZN(p7_S[63]) );
  XNOR2_X1 U971 ( .A(n879), .B(n858), .ZN(n714) );
  XNOR2_X1 U999 ( .A(n880), .B(n881), .ZN(n900) );
  AOI22_X1 U1035 ( .A1(B1[4]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_17_), .ZN(n923) );
  OAI221_X1 U1034 ( .B1(B1[3]), .B2(n763), .C1(p7_minus_A_shifted_16_), .C2(
        n764), .A(n923), .ZN(n913) );
  AOI222_X1 U1021 ( .A1(p7_muxs_out_2__12_), .A2(p7_muxs_out_3__12_), .B1(
        p7_muxs_out_2__12_), .B2(n913), .C1(p7_muxs_out_3__12_), .C2(n913), 
        .ZN(n873) );
  AOI22_X1 U1015 ( .A1(B1[0]), .A2(n668), .B1(n667), .B2(
        p7_minus_A_shifted_13_), .ZN(n909) );
  AOI221_X1 U1014 ( .B1(n670), .B2(B1[1]), .C1(n671), .C2(
        p7_minus_A_shifted_14_), .A(n909), .ZN(n874) );
  XNOR2_X1 U1013 ( .A(n873), .B(n874), .ZN(n907) );
  AOI22_X1 U1012 ( .A1(B1[3]), .A2(n751), .B1(n752), .B2(
        p7_minus_A_shifted_16_), .ZN(n908) );
  OAI221_X1 U1011 ( .B1(B1[2]), .B2(n748), .C1(p7_minus_A_shifted_15_), .C2(
        n749), .A(n908), .ZN(n875) );
  XNOR2_X1 U1010 ( .A(n907), .B(n875), .ZN(n877) );
  XNOR2_X1 U1032 ( .A(p7_muxs_out_2__12_), .B(n922), .ZN(n897) );
  OAI21_X1 U1028 ( .B1(n919), .B2(p7_muxs_out_1__12_), .A(n882), .ZN(n898) );
  AOI22_X1 U1054 ( .A1(n943), .A2(p7_minus_A_shifted_23_), .B1(n886), .B2(
        B1[11]), .ZN(n942) );
  OAI21_X1 U1053 ( .B1(B1[11]), .B2(n920), .A(n942), .ZN(n941) );
  NAND2_X1 U1052 ( .A1(p7_muxs_out_1__11_), .A2(n941), .ZN(n899) );
  AOI222_X1 U996 ( .A1(n897), .A2(n898), .B1(n897), .B2(n899), .C1(n898), .C2(
        n899), .ZN(n878) );
  AOI222_X1 U970 ( .A1(n876), .A2(n877), .B1(n876), .B2(n878), .C1(n877), .C2(
        n878), .ZN(n715) );
  OAI222_X1 U968 ( .A1(n872), .A2(n873), .B1(n872), .B2(n874), .C1(n873), .C2(
        n874), .ZN(n871) );
  AOI222_X1 U966 ( .A1(n714), .A2(n715), .B1(n714), .B2(n712), .C1(n715), .C2(
        n712), .ZN(p7_C[62]) );
  XNOR2_X1 U803 ( .A(n712), .B(n713), .ZN(p7_S[62]) );
  XNOR2_X1 U995 ( .A(n896), .B(n878), .ZN(n718) );
  AOI22_X1 U1041 ( .A1(B1[2]), .A2(n751), .B1(n752), .B2(
        p7_minus_A_shifted_15_), .ZN(n927) );
  OAI221_X1 U1040 ( .B1(B1[1]), .B2(n748), .C1(p7_minus_A_shifted_14_), .C2(
        n749), .A(n927), .ZN(n891) );
  NOR2_X1 U1038 ( .A1(n910), .A2(p7_minus_A_shifted_13_), .ZN(n924) );
  XNOR2_X1 U1027 ( .A(n897), .B(n898), .ZN(n918) );
  OAI21_X1 U1051 ( .B1(p7_muxs_out_1__11_), .B2(n941), .A(n899), .ZN(n928) );
  AOI22_X1 U1078 ( .A1(n943), .A2(p7_minus_A_shifted_22_), .B1(n886), .B2(
        B1[10]), .ZN(n956) );
  OAI21_X1 U1077 ( .B1(B1[10]), .B2(n920), .A(n956), .ZN(n955) );
  NAND2_X1 U1076 ( .A1(p7_muxs_out_1__10_), .A2(n955), .ZN(n930) );
  AOI222_X1 U1042 ( .A1(n928), .A2(n929), .B1(n928), .B2(n930), .C1(n929), 
        .C2(n930), .ZN(n895) );
  AOI222_X1 U994 ( .A1(n893), .A2(n894), .B1(n893), .B2(n895), .C1(n894), .C2(
        n895), .ZN(n719) );
  OAI221_X1 U991 ( .B1(B1[0]), .B2(n756), .C1(p7_minus_A_shifted_13_), .C2(
        n755), .A(n667), .ZN(n892) );
  AOI222_X1 U990 ( .A1(n891), .A2(reg2_reg[13]), .B1(n891), .B2(n892), .C1(
        reg2_reg[13]), .C2(n892), .ZN(n716) );
  AOI222_X1 U989 ( .A1(n718), .A2(n719), .B1(n718), .B2(n716), .C1(n719), .C2(
        n716), .ZN(p7_C[61]) );
  XNOR2_X1 U805 ( .A(n716), .B(n717), .ZN(p7_S[61]) );
  AOI22_X1 U1065 ( .A1(B1[1]), .A2(n751), .B1(n752), .B2(
        p7_minus_A_shifted_14_), .ZN(n947) );
  OAI221_X1 U1064 ( .B1(B1[0]), .B2(n748), .C1(p7_minus_A_shifted_13_), .C2(
        n749), .A(n947), .ZN(n931) );
  AOI22_X1 U1061 ( .A1(B1[3]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_16_), .ZN(n946) );
  OAI221_X1 U1060 ( .B1(B1[2]), .B2(n763), .C1(p7_minus_A_shifted_15_), .C2(
        n764), .A(n946), .ZN(n932) );
  AOI222_X1 U1043 ( .A1(n931), .A2(p7_muxs_out_3__11_), .B1(n931), .B2(n932), 
        .C1(p7_muxs_out_3__11_), .C2(n932), .ZN(n722) );
  XNOR2_X1 U1024 ( .A(n895), .B(n917), .ZN(n723) );
  XNOR2_X1 U1063 ( .A(n931), .B(p7_muxs_out_3__11_), .ZN(n945) );
  XNOR2_X1 U1059 ( .A(n945), .B(n932), .ZN(n914) );
  AOI22_X1 U1056 ( .A1(p7_muxs_out_2__11_), .A2(n944), .B1(n930), .B2(n929), 
        .ZN(n940) );
  XNOR2_X1 U1050 ( .A(n940), .B(n928), .ZN(n915) );
  OAI21_X1 U1075 ( .B1(p7_muxs_out_1__10_), .B2(n955), .A(n930), .ZN(n951) );
  AOI222_X1 U1069 ( .A1(n949), .A2(n950), .B1(n949), .B2(n951), .C1(n950), 
        .C2(n951), .ZN(n916) );
  AOI222_X1 U1023 ( .A1(n914), .A2(n915), .B1(n914), .B2(n916), .C1(n915), 
        .C2(n916), .ZN(n720) );
  AOI222_X1 U1022 ( .A1(n722), .A2(n723), .B1(n722), .B2(n720), .C1(n723), 
        .C2(n720), .ZN(p7_C[60]) );
  AOI22_X1 U1087 ( .A1(B1[2]), .A2(n772), .B1(n773), .B2(
        p7_minus_A_shifted_15_), .ZN(n957) );
  OAI221_X1 U1086 ( .B1(B1[1]), .B2(n763), .C1(p7_minus_A_shifted_14_), .C2(
        n764), .A(n957), .ZN(n934) );
  NOR2_X1 U1083 ( .A1(n948), .A2(p7_minus_A_shifted_13_), .ZN(n935) );
  XNOR2_X1 U1048 ( .A(n916), .B(n939), .ZN(n726) );
  AOI22_X1 U1079 ( .A1(p7_muxs_out_2__10_), .A2(p7_muxs_out_3__10_), .B1(n950), 
        .B2(n949), .ZN(n954) );
  XNOR2_X1 U1074 ( .A(n954), .B(n951), .ZN(n937) );
  NOR2_X1 U1103 ( .A1(B1[8]), .A2(n902), .ZN(n972) );
  AOI221_X1 U1102 ( .B1(B1[9]), .B2(n886), .C1(p7_minus_A_shifted_22_), .C2(
        n904), .A(n972), .ZN(n960) );
  AOI222_X1 U1089 ( .A1(n958), .A2(n959), .B1(n958), .B2(n960), .C1(n959), 
        .C2(n960), .ZN(n938) );
  AOI222_X1 U1047 ( .A1(n936), .A2(n937), .B1(n936), .B2(n938), .C1(n937), 
        .C2(n938), .ZN(n727) );
  AOI22_X1 U1105 ( .A1(p7_muxs_out_1__9_), .A2(p7_muxs_out_2__9_), .B1(n959), 
        .B2(n958), .ZN(n971) );
  XNOR2_X1 U1101 ( .A(n971), .B(n960), .ZN(n961) );
  AOI22_X1 U1099 ( .A1(B1[0]), .A2(n764), .B1(n763), .B2(
        p7_minus_A_shifted_13_), .ZN(n970) );
  OAI221_X1 U1097 ( .B1(n967), .B2(p7_minus_A_shifted_14_), .C1(n968), .C2(
        B1[1]), .A(n969), .ZN(n952) );
  AOI22_X1 U1126 ( .A1(B1[8]), .A2(n886), .B1(n904), .B2(
        p7_minus_A_shifted_21_), .ZN(n982) );
  OAI21_X1 U1125 ( .B1(B1[7]), .B2(n902), .A(n982), .ZN(n966) );
  AOI222_X1 U1094 ( .A1(p7_muxs_out_1__8_), .A2(p7_muxs_out_2__8_), .B1(
        p7_muxs_out_1__8_), .B2(n966), .C1(p7_muxs_out_2__8_), .C2(n966), .ZN(
        n964) );
  AOI222_X1 U1090 ( .A1(n961), .A2(n962), .B1(n961), .B2(n963), .C1(n962), 
        .C2(n963), .ZN(n730) );
  XNOR2_X1 U1072 ( .A(n938), .B(n953), .ZN(n731) );
  NAND2_X1 U1071 ( .A1(p7_muxs_out_3__9_), .A2(n952), .ZN(n728) );
  XNOR2_X1 U1095 ( .A(n961), .B(n962), .ZN(n965) );
  XNOR2_X1 U1093 ( .A(n965), .B(n964), .ZN(n732) );
  OAI221_X1 U1115 ( .B1(n967), .B2(p7_minus_A_shifted_13_), .C1(n968), .C2(
        B1[0]), .A(n763), .ZN(n973) );
  AOI22_X1 U1139 ( .A1(B1[7]), .A2(n921), .B1(n920), .B2(
        p7_minus_A_shifted_20_), .ZN(n988) );
  AOI21_X1 U1138 ( .B1(n943), .B2(p7_minus_A_shifted_19_), .A(n988), .ZN(n986)
         );
  NOR2_X1 U1136 ( .A1(n986), .A2(n2855), .ZN(n975) );
  XNOR2_X1 U1128 ( .A(p7_muxs_out_2__8_), .B(p7_muxs_out_1__8_), .ZN(n981) );
  XNOR2_X1 U1124 ( .A(n981), .B(n966), .ZN(n976) );
  AOI222_X1 U1109 ( .A1(n974), .A2(n975), .B1(n974), .B2(n976), .C1(n975), 
        .C2(n976), .ZN(n734) );
  NAND2_X1 U1108 ( .A1(p7_muxs_out_3__8_), .A2(n973), .ZN(n735) );
  XNOR2_X1 U1112 ( .A(n976), .B(n979), .ZN(n736) );
  NOR2_X1 U1148 ( .A1(B1[5]), .A2(n902), .ZN(n991) );
  AOI221_X1 U1147 ( .B1(B1[6]), .B2(n886), .C1(p7_minus_A_shifted_19_), .C2(
        n904), .A(n991), .ZN(n984) );
  NOR2_X1 U1133 ( .A1(n984), .A2(n985), .ZN(n977) );
  AOI22_X1 U816 ( .A1(reg2_reg[9]), .A2(n738), .B1(n739), .B2(n2812), .ZN(n737) );
  XNOR2_X1 U815 ( .A(n736), .B(n737), .ZN(p7_S[56]) );
  XNOR2_X1 U1146 ( .A(p7_muxs_out_1__6_), .B(n984), .ZN(n990) );
  NAND2_X1 U1145 ( .A1(n990), .A2(p7_muxs_out_2__6_), .ZN(n744) );
  AOI222_X1 U1129 ( .A1(n742), .A2(n745), .B1(n742), .B2(n744), .C1(n745), 
        .C2(n744), .ZN(p7_C[55]) );
  AOI22_X1 U819 ( .A1(p7_muxs_out_3__7_), .A2(n743), .B1(n744), .B2(n745), 
        .ZN(n741) );
  XNOR2_X1 U818 ( .A(n741), .B(n742), .ZN(p7_S[55]) );
  OAI21_X1 U1144 ( .B1(n990), .B2(p7_muxs_out_2__6_), .A(n744), .ZN(n746) );
  NOR2_X1 U1143 ( .A1(n989), .A2(n746), .ZN(p7_C[54]) );
  XNOR2_X1 U821 ( .A(p7_muxs_out_3__6_), .B(n746), .ZN(p7_S[54]) );
  AOI222_X1 U1044 ( .A1(n726), .A2(n727), .B1(n726), .B2(n724), .C1(n727), 
        .C2(n724), .ZN(p7_C[59]) );
  XNOR2_X1 U807 ( .A(n720), .B(n721), .ZN(p7_S[60]) );
  NAND2_X1 U2420 ( .A1(VIN), .A2(temp1[12]), .ZN(n2059) );
  OAI21_X1 U2419 ( .B1(VIN), .B2(n2187), .A(n2059), .ZN(n2448) );
  NAND2_X1 U2356 ( .A1(VIN), .A2(temp3[12]), .ZN(n2029) );
  OAI21_X1 U2355 ( .B1(VIN), .B2(n2158), .A(n2029), .ZN(n2416) );
  NAND2_X1 U2388 ( .A1(VIN), .A2(temp2[12]), .ZN(n2044) );
  OAI21_X1 U2387 ( .B1(VIN), .B2(n2173), .A(n2044), .ZN(n2432) );
  NAND2_X1 U2322 ( .A1(VIN), .A2(temp4[12]), .ZN(n2013) );
  OAI21_X1 U2321 ( .B1(VIN), .B2(n2143), .A(n2013), .ZN(n2399) );
  NAND2_X1 U2422 ( .A1(VIN), .A2(temp1[11]), .ZN(n2060) );
  OAI21_X1 U2421 ( .B1(VIN), .B2(n2188), .A(n2060), .ZN(n2449) );
  NAND2_X1 U2324 ( .A1(VIN), .A2(temp4[11]), .ZN(n2014) );
  OAI21_X1 U2323 ( .B1(VIN), .B2(n2144), .A(n2014), .ZN(n2400) );
  NAND2_X1 U2390 ( .A1(VIN), .A2(temp2[11]), .ZN(n2045) );
  OAI21_X1 U2389 ( .B1(VIN), .B2(n2174), .A(n2045), .ZN(n2433) );
  NAND2_X1 U2358 ( .A1(VIN), .A2(temp3[11]), .ZN(n2030) );
  OAI21_X1 U2357 ( .B1(VIN), .B2(n2159), .A(n2030), .ZN(n2417) );
  NAND2_X1 U2424 ( .A1(VIN), .A2(temp1[10]), .ZN(n2061) );
  OAI21_X1 U2423 ( .B1(VIN), .B2(n2189), .A(n2061), .ZN(n2450) );
  NAND2_X1 U2392 ( .A1(VIN), .A2(temp2[10]), .ZN(n2046) );
  OAI21_X1 U2391 ( .B1(VIN), .B2(n2175), .A(n2046), .ZN(n2434) );
  NAND2_X1 U2360 ( .A1(VIN), .A2(temp3[10]), .ZN(n2031) );
  OAI21_X1 U2359 ( .B1(VIN), .B2(n2160), .A(n2031), .ZN(n2418) );
  NAND2_X1 U2326 ( .A1(VIN), .A2(temp4[10]), .ZN(n2015) );
  OAI21_X1 U2325 ( .B1(VIN), .B2(n2145), .A(n2015), .ZN(n2401) );
  NAND2_X1 U2426 ( .A1(VIN), .A2(temp1[9]), .ZN(n2062) );
  OAI21_X1 U2425 ( .B1(VIN), .B2(n2190), .A(n2062), .ZN(n2451) );
  NAND2_X1 U2328 ( .A1(VIN), .A2(temp4[9]), .ZN(n2016) );
  OAI21_X1 U2327 ( .B1(VIN), .B2(n2146), .A(n2016), .ZN(n2402) );
  NAND2_X1 U2394 ( .A1(VIN), .A2(temp2[9]), .ZN(n2047) );
  OAI21_X1 U2393 ( .B1(VIN), .B2(n2176), .A(n2047), .ZN(n2435) );
  NAND2_X1 U2362 ( .A1(VIN), .A2(temp3[9]), .ZN(n2032) );
  OAI21_X1 U2361 ( .B1(VIN), .B2(n2161), .A(n2032), .ZN(n2419) );
  NAND2_X1 U2428 ( .A1(VIN), .A2(temp1[8]), .ZN(n2063) );
  OAI21_X1 U2427 ( .B1(VIN), .B2(n2191), .A(n2063), .ZN(n2452) );
  NAND2_X1 U2364 ( .A1(VIN), .A2(temp3[8]), .ZN(n2033) );
  OAI21_X1 U2363 ( .B1(VIN), .B2(n2162), .A(n2033), .ZN(n2420) );
  NAND2_X1 U2330 ( .A1(VIN), .A2(temp4[8]), .ZN(n2017) );
  OAI21_X1 U2329 ( .B1(VIN), .B2(n2147), .A(n2017), .ZN(n2403) );
  NAND2_X1 U2396 ( .A1(VIN), .A2(temp2[8]), .ZN(n2048) );
  OAI21_X1 U2395 ( .B1(VIN), .B2(n2177), .A(n2048), .ZN(n2436) );
  NAND2_X1 U2430 ( .A1(VIN), .A2(temp1[7]), .ZN(n2064) );
  OAI21_X1 U2429 ( .B1(VIN), .B2(n2192), .A(n2064), .ZN(n2453) );
  NAND2_X1 U2366 ( .A1(VIN), .A2(temp3[7]), .ZN(n2034) );
  OAI21_X1 U2365 ( .B1(VIN), .B2(n2163), .A(n2034), .ZN(n2421) );
  NAND2_X1 U2332 ( .A1(VIN), .A2(temp4[7]), .ZN(n2018) );
  OAI21_X1 U2331 ( .B1(VIN), .B2(n2148), .A(n2018), .ZN(n2404) );
  NAND2_X1 U2398 ( .A1(VIN), .A2(temp2[7]), .ZN(n2049) );
  OAI21_X1 U2397 ( .B1(VIN), .B2(n2178), .A(n2049), .ZN(n2437) );
  NAND2_X1 U2432 ( .A1(VIN), .A2(temp1[6]), .ZN(n2065) );
  OAI21_X1 U2431 ( .B1(VIN), .B2(n2193), .A(n2065), .ZN(n2454) );
  NAND2_X1 U2368 ( .A1(VIN), .A2(temp3[6]), .ZN(n2035) );
  OAI21_X1 U2367 ( .B1(VIN), .B2(n2164), .A(n2035), .ZN(n2422) );
  NAND2_X1 U2400 ( .A1(VIN), .A2(temp2[6]), .ZN(n2050) );
  OAI21_X1 U2399 ( .B1(VIN), .B2(n2179), .A(n2050), .ZN(n2438) );
  NAND2_X1 U2334 ( .A1(VIN), .A2(temp4[6]), .ZN(n2019) );
  OAI21_X1 U2333 ( .B1(VIN), .B2(n2149), .A(n2019), .ZN(n2405) );
  NAND2_X1 U2434 ( .A1(VIN), .A2(temp1[5]), .ZN(n2066) );
  OAI21_X1 U2433 ( .B1(VIN), .B2(n2194), .A(n2066), .ZN(n2455) );
  NAND2_X1 U2402 ( .A1(VIN), .A2(temp2[5]), .ZN(n2051) );
  OAI21_X1 U2401 ( .B1(VIN), .B2(n2180), .A(n2051), .ZN(n2439) );
  NAND2_X1 U2370 ( .A1(VIN), .A2(temp3[5]), .ZN(n2036) );
  OAI21_X1 U2369 ( .B1(VIN), .B2(n2165), .A(n2036), .ZN(n2423) );
  NAND2_X1 U2336 ( .A1(VIN), .A2(temp4[5]), .ZN(n2020) );
  OAI21_X1 U2335 ( .B1(VIN), .B2(n2150), .A(n2020), .ZN(n2406) );
  NAND2_X1 U2436 ( .A1(VIN), .A2(temp1[4]), .ZN(n2067) );
  OAI21_X1 U2435 ( .B1(VIN), .B2(n2195), .A(n2067), .ZN(n2456) );
  NAND2_X1 U2372 ( .A1(VIN), .A2(temp3[4]), .ZN(n2037) );
  OAI21_X1 U2371 ( .B1(VIN), .B2(n2166), .A(n2037), .ZN(n2424) );
  NAND2_X1 U2404 ( .A1(VIN), .A2(temp2[4]), .ZN(n2052) );
  OAI21_X1 U2403 ( .B1(VIN), .B2(n2181), .A(n2052), .ZN(n2440) );
  NAND2_X1 U2338 ( .A1(VIN), .A2(temp4[4]), .ZN(n2021) );
  OAI21_X1 U2337 ( .B1(VIN), .B2(n2151), .A(n2021), .ZN(n2407) );
  NAND2_X1 U2438 ( .A1(VIN), .A2(temp1[3]), .ZN(n2068) );
  OAI21_X1 U2437 ( .B1(VIN), .B2(n2196), .A(n2068), .ZN(n2457) );
  NAND2_X1 U2406 ( .A1(VIN), .A2(temp2[3]), .ZN(n2053) );
  OAI21_X1 U2405 ( .B1(VIN), .B2(n2182), .A(n2053), .ZN(n2441) );
  NAND2_X1 U2340 ( .A1(VIN), .A2(temp4[3]), .ZN(n2022) );
  OAI21_X1 U2339 ( .B1(VIN), .B2(n2152), .A(n2022), .ZN(n2408) );
  NAND2_X1 U2374 ( .A1(VIN), .A2(temp3[3]), .ZN(n2038) );
  OAI21_X1 U2373 ( .B1(VIN), .B2(n2167), .A(n2038), .ZN(n2425) );
  NAND2_X1 U2440 ( .A1(VIN), .A2(temp1[2]), .ZN(n2069) );
  OAI21_X1 U2439 ( .B1(VIN), .B2(n2197), .A(n2069), .ZN(n2458) );
  NAND2_X1 U2408 ( .A1(VIN), .A2(temp2[2]), .ZN(n2054) );
  OAI21_X1 U2407 ( .B1(VIN), .B2(n2183), .A(n2054), .ZN(n2442) );
  NAND2_X1 U2342 ( .A1(VIN), .A2(temp4[2]), .ZN(n2023) );
  OAI21_X1 U2341 ( .B1(VIN), .B2(n2153), .A(n2023), .ZN(n2409) );
  NAND2_X1 U2376 ( .A1(VIN), .A2(temp3[2]), .ZN(n2039) );
  OAI21_X1 U2375 ( .B1(VIN), .B2(n2168), .A(n2039), .ZN(n2426) );
  NAND2_X1 U2442 ( .A1(VIN), .A2(temp1[1]), .ZN(n2070) );
  OAI21_X1 U2441 ( .B1(VIN), .B2(n2198), .A(n2070), .ZN(n2459) );
  NAND2_X1 U2344 ( .A1(VIN), .A2(temp4[1]), .ZN(n2024) );
  OAI21_X1 U2343 ( .B1(VIN), .B2(n2154), .A(n2024), .ZN(n2410) );
  NAND2_X1 U2378 ( .A1(VIN), .A2(temp3[1]), .ZN(n2040) );
  OAI21_X1 U2377 ( .B1(VIN), .B2(n2169), .A(n2040), .ZN(n2427) );
  NAND2_X1 U2410 ( .A1(VIN), .A2(temp2[1]), .ZN(n2055) );
  OAI21_X1 U2409 ( .B1(VIN), .B2(n2184), .A(n2055), .ZN(n2443) );
  NAND2_X1 U2444 ( .A1(VIN), .A2(temp1[0]), .ZN(n2071) );
  OAI21_X1 U2443 ( .B1(VIN), .B2(n2199), .A(n2071), .ZN(n2460) );
  NAND2_X1 U2412 ( .A1(VIN), .A2(temp2[0]), .ZN(n2056) );
  OAI21_X1 U2411 ( .B1(VIN), .B2(n2185), .A(n2056), .ZN(n2444) );
  NAND2_X1 U2380 ( .A1(VIN), .A2(temp3[0]), .ZN(n2041) );
  OAI21_X1 U2379 ( .B1(VIN), .B2(n2170), .A(n2041), .ZN(n2428) );
  NAND2_X1 U2346 ( .A1(VIN), .A2(temp4[0]), .ZN(n2025) );
  OAI21_X1 U2345 ( .B1(VIN), .B2(n2155), .A(n2025), .ZN(n2411) );
  OAI21_X1 U2415 ( .B1(VIN), .B2(n2860), .A(n2057), .ZN(n2446) );
  OAI21_X1 U2445 ( .B1(VIN), .B2(n2867), .A(n2057), .ZN(n2461) );
  NAND2_X1 U2292 ( .A1(VIN), .A2(ff[13]), .ZN(n1998) );
  OAI21_X1 U2291 ( .B1(VIN), .B2(n2128), .A(n1998), .ZN(n2384) );
  NAND2_X1 U2294 ( .A1(VIN), .A2(ff[12]), .ZN(n1999) );
  OAI21_X1 U2293 ( .B1(VIN), .B2(n2129), .A(n1999), .ZN(n2385) );
  NAND2_X1 U2463 ( .A1(VIN), .A2(w[12]), .ZN(n2074) );
  OAI21_X1 U2460 ( .B1(VIN), .B2(n2863), .A(n2074), .ZN(n2468) );
  OAI21_X1 U2462 ( .B1(VIN), .B2(n2848), .A(n2074), .ZN(n2469) );
  NAND2_X1 U2296 ( .A1(VIN), .A2(ff[11]), .ZN(n2000) );
  OAI21_X1 U2295 ( .B1(VIN), .B2(n2130), .A(n2000), .ZN(n2386) );
  NAND2_X1 U2480 ( .A1(VIN), .A2(w[11]), .ZN(n2077) );
  OAI21_X1 U2477 ( .B1(VIN), .B2(n2862), .A(n2077), .ZN(n2476) );
  OAI21_X1 U2479 ( .B1(VIN), .B2(n2790), .A(n2077), .ZN(n2477) );
  NAND2_X1 U2298 ( .A1(VIN), .A2(ff[10]), .ZN(n2001) );
  OAI21_X1 U2297 ( .B1(VIN), .B2(n2131), .A(n2001), .ZN(n2387) );
  NAND2_X1 U2497 ( .A1(VIN), .A2(w[10]), .ZN(n2083) );
  OAI21_X1 U2494 ( .B1(VIN), .B2(n2833), .A(n2083), .ZN(n2484) );
  OAI21_X1 U2496 ( .B1(VIN), .B2(n2880), .A(n2083), .ZN(n2485) );
  NAND2_X1 U2300 ( .A1(VIN), .A2(ff[9]), .ZN(n2002) );
  OAI21_X1 U2299 ( .B1(VIN), .B2(n2132), .A(n2002), .ZN(n2388) );
  NAND2_X1 U2514 ( .A1(VIN), .A2(w[9]), .ZN(n2087) );
  OAI21_X1 U2511 ( .B1(VIN), .B2(n2816), .A(n2087), .ZN(n2492) );
  OAI21_X1 U2513 ( .B1(VIN), .B2(n2819), .A(n2087), .ZN(n2493) );
  NAND2_X1 U2302 ( .A1(VIN), .A2(ff[8]), .ZN(n2003) );
  OAI21_X1 U2301 ( .B1(VIN), .B2(n2133), .A(n2003), .ZN(n2389) );
  NAND2_X1 U2531 ( .A1(VIN), .A2(w[8]), .ZN(n2093) );
  OAI21_X1 U2528 ( .B1(VIN), .B2(n2811), .A(n2093), .ZN(n2500) );
  OAI21_X1 U2530 ( .B1(VIN), .B2(n2881), .A(n2093), .ZN(n2501) );
  NAND2_X1 U2304 ( .A1(VIN), .A2(ff[7]), .ZN(n2004) );
  OAI21_X1 U2303 ( .B1(VIN), .B2(n2134), .A(n2004), .ZN(n2390) );
  NAND2_X1 U2548 ( .A1(VIN), .A2(w[7]), .ZN(n2100) );
  OAI21_X1 U2545 ( .B1(VIN), .B2(n2831), .A(n2100), .ZN(n2508) );
  OAI21_X1 U2547 ( .B1(VIN), .B2(n2796), .A(n2100), .ZN(n2509) );
  NAND2_X1 U2306 ( .A1(VIN), .A2(ff[6]), .ZN(n2005) );
  OAI21_X1 U2305 ( .B1(VIN), .B2(n2135), .A(n2005), .ZN(n2391) );
  NAND2_X1 U2560 ( .A1(VIN), .A2(w[6]), .ZN(n2104) );
  OAI21_X1 U2559 ( .B1(VIN), .B2(n2835), .A(n2104), .ZN(n2516) );
  NAND2_X1 U2308 ( .A1(VIN), .A2(ff[5]), .ZN(n2006) );
  OAI21_X1 U2307 ( .B1(VIN), .B2(n2136), .A(n2006), .ZN(n2392) );
  NAND2_X1 U2573 ( .A1(VIN), .A2(w[5]), .ZN(n2107) );
  OAI21_X1 U2572 ( .B1(VIN), .B2(n2834), .A(n2107), .ZN(n2524) );
  AOI22_X1 U2553 ( .A1(VIN), .A2(n2835), .B1(n2815), .B2(n3435), .ZN(n2512) );
  AOI22_X1 U2503 ( .A1(VIN), .A2(n2816), .B1(n2814), .B2(n3435), .ZN(n2488) );
  AOI22_X1 U2413 ( .A1(VIN), .A2(n2860), .B1(n2866), .B2(n3435), .ZN(n2445) );
  AOI22_X1 U2383 ( .A1(VIN), .A2(n2860), .B1(n2878), .B2(n3435), .ZN(n2430) );
  AOI22_X1 U2452 ( .A1(VIN), .A2(n2863), .B1(n2858), .B2(n3435), .ZN(n2464) );
  AOI22_X1 U2537 ( .A1(VIN), .A2(n2831), .B1(n2830), .B2(n3435), .ZN(n2504) );
  AOI22_X1 U2556 ( .A1(VIN), .A2(n2835), .B1(n2896), .B2(n3435), .ZN(n2514) );
  AOI22_X1 U2509 ( .A1(VIN), .A2(n2816), .B1(n2812), .B2(n3435), .ZN(n2491) );
  AOI22_X1 U2507 ( .A1(VIN), .A2(n2816), .B1(n2872), .B2(n3435), .ZN(n2490) );
  AOI22_X1 U2543 ( .A1(VIN), .A2(n2831), .B1(n2799), .B2(n3435), .ZN(n2507) );
  AOI22_X1 U2458 ( .A1(VIN), .A2(n2863), .B1(n2849), .B2(n3435), .ZN(n2467) );
  AOI22_X1 U2456 ( .A1(VIN), .A2(n2863), .B1(n2876), .B2(n3435), .ZN(n2466) );
  AOI22_X1 U2541 ( .A1(VIN), .A2(n2831), .B1(n2870), .B2(n3435), .ZN(n2506) );
  AOI22_X1 U2524 ( .A1(VIN), .A2(n2811), .B1(n2806), .B2(n3435), .ZN(n2498) );
  AOI22_X1 U2492 ( .A1(VIN), .A2(n2833), .B1(n2882), .B2(n3435), .ZN(n2483) );
  AOI22_X1 U2526 ( .A1(VIN), .A2(n2811), .B1(n2885), .B2(n3435), .ZN(n2499) );
  AOI22_X1 U2486 ( .A1(VIN), .A2(n2833), .B1(n2810), .B2(n3435), .ZN(n2480) );
  AOI22_X1 U2551 ( .A1(VIN), .A2(n2815), .B1(n2897), .B2(n3435), .ZN(n2511) );
  AOI22_X1 U2490 ( .A1(VIN), .A2(n2833), .B1(n2808), .B2(n3435), .ZN(n2482) );
  AOI22_X1 U2520 ( .A1(VIN), .A2(n2811), .B1(n2832), .B2(n3435), .ZN(n2496) );
  AOI22_X1 U2475 ( .A1(VIN), .A2(n2862), .B1(n2791), .B2(n3435), .ZN(n2475) );
  AOI22_X1 U2469 ( .A1(VIN), .A2(n2862), .B1(n2861), .B2(n3435), .ZN(n2472) );
  AOI22_X1 U2473 ( .A1(VIN), .A2(n2862), .B1(n2874), .B2(n3435), .ZN(n2474) );
  AOI22_X1 U2450 ( .A1(VIN), .A2(n2858), .B1(n2877), .B2(n3435), .ZN(n2463) );
  AOI22_X1 U2501 ( .A1(VIN), .A2(n2814), .B1(n2873), .B2(n3435), .ZN(n2487) );
  AOI22_X1 U2535 ( .A1(VIN), .A2(n2830), .B1(n2871), .B2(n3435), .ZN(n2503) );
  AOI22_X1 U2569 ( .A1(VIN), .A2(n2834), .B1(n2894), .B2(n3435), .ZN(n2522) );
  AOI22_X1 U2582 ( .A1(VIN), .A2(n2817), .B1(n2892), .B2(n3435), .ZN(n2530) );
  AOI22_X1 U2518 ( .A1(VIN), .A2(n2832), .B1(n2807), .B2(n3435), .ZN(n2495) );
  AOI22_X1 U2579 ( .A1(VIN), .A2(n2817), .B1(n2818), .B2(n3435), .ZN(n2528) );
  AOI22_X1 U2484 ( .A1(VIN), .A2(n2810), .B1(n2809), .B2(n3435), .ZN(n2479) );
  AOI22_X1 U2566 ( .A1(VIN), .A2(n2834), .B1(n2813), .B2(n3435), .ZN(n2520) );
  AOI22_X1 U2467 ( .A1(VIN), .A2(n2861), .B1(n2875), .B2(n3435), .ZN(n2471) );
  AOI22_X1 U2577 ( .A1(VIN), .A2(n2818), .B1(n2893), .B2(n3435), .ZN(n2527) );
  AOI22_X1 U2592 ( .A1(VIN), .A2(p11_minus_A_shifted_16_), .B1(
        p10_minus_A_shifted_16_), .B2(n3435), .ZN(n2536) );
  AOI22_X1 U2564 ( .A1(VIN), .A2(n2813), .B1(n2895), .B2(n3435), .ZN(n2519) );
  AOI22_X1 U2595 ( .A1(VIN), .A2(p11_minus_A_shifted_16_), .B1(n2890), .B2(
        n3435), .ZN(n2538) );
  AOI22_X1 U2625 ( .A1(VIN), .A2(p11_minus_A_shifted_14_), .B1(n2865), .B2(
        n3435), .ZN(n2555) );
  AOI22_X1 U2605 ( .A1(VIN), .A2(n2820), .B1(n2821), .B2(n3435), .ZN(n2544) );
  AOI22_X1 U2608 ( .A1(VIN), .A2(n2820), .B1(n2888), .B2(n3435), .ZN(n2546) );
  AOI22_X1 U2619 ( .A1(VIN), .A2(p11_minus_A_shifted_14_), .B1(
        p10_minus_A_shifted_14_), .B2(n3435), .ZN(n2552) );
  AOI22_X1 U2590 ( .A1(VIN), .A2(p10_minus_A_shifted_16_), .B1(n2891), .B2(
        n3435), .ZN(n2535) );
  AOI22_X1 U2603 ( .A1(VIN), .A2(n2821), .B1(n2889), .B2(n3435), .ZN(n2543) );
  AOI22_X1 U2634 ( .A1(VIN), .A2(n2839), .B1(n2869), .B2(n3435), .ZN(n2559) );
  AOI22_X1 U2638 ( .A1(VIN), .A2(n2868), .B1(n2797), .B2(n3435), .ZN(n2561) );
  AOI22_X1 U2632 ( .A1(VIN), .A2(n2869), .B1(n2798), .B2(n3435), .ZN(n2558) );
  AOI22_X1 U2499 ( .A1(VIN), .A2(n2873), .B1(n2789), .B2(n3435), .ZN(n2486) );
  AOI22_X1 U2482 ( .A1(VIN), .A2(n2809), .B1(n2884), .B2(n3435), .ZN(n2478) );
  AOI22_X1 U2448 ( .A1(VIN), .A2(n2877), .B1(n2803), .B2(n3435), .ZN(n2462) );
  AOI22_X1 U2454 ( .A1(VIN), .A2(n2876), .B1(n2802), .B2(n3435), .ZN(n2465) );
  AOI22_X1 U2465 ( .A1(VIN), .A2(n2875), .B1(n2787), .B2(n3435), .ZN(n2470) );
  AOI22_X1 U2471 ( .A1(VIN), .A2(n2874), .B1(n2786), .B2(n3435), .ZN(n2473) );
  AOI22_X1 U2381 ( .A1(VIN), .A2(n2878), .B1(n2805), .B2(n3435), .ZN(n2429) );
  AOI22_X1 U2539 ( .A1(VIN), .A2(n2870), .B1(n2800), .B2(n3435), .ZN(n2505) );
  AOI22_X1 U2522 ( .A1(VIN), .A2(n2806), .B1(n2886), .B2(n3435), .ZN(n2497) );
  AOI22_X1 U2488 ( .A1(VIN), .A2(n2808), .B1(n2883), .B2(n3435), .ZN(n2481) );
  AOI22_X1 U2533 ( .A1(VIN), .A2(n2871), .B1(n2801), .B2(n3435), .ZN(n2502) );
  AOI22_X1 U2505 ( .A1(VIN), .A2(n2872), .B1(n2788), .B2(n3435), .ZN(n2489) );
  AOI22_X1 U2516 ( .A1(VIN), .A2(n2807), .B1(n2887), .B2(n3435), .ZN(n2494) );
  NAND2_X1 U2665 ( .A1(n2226), .A2(n3435), .ZN(n2581) );
  NAND2_X1 U2310 ( .A1(VIN), .A2(ff[4]), .ZN(n2007) );
  OAI21_X1 U2309 ( .B1(VIN), .B2(n2137), .A(n2007), .ZN(n2393) );
  NAND2_X1 U2586 ( .A1(VIN), .A2(w[4]), .ZN(n2110) );
  OAI21_X1 U2585 ( .B1(VIN), .B2(n2817), .A(n2110), .ZN(n2532) );
  OAI22_X1 U2618 ( .A1(n3435), .A2(reg4[1]), .B1(n2222), .B2(VIN), .ZN(n2118)
         );
  OAI22_X1 U2624 ( .A1(n3435), .A2(reg2[1]), .B1(n2223), .B2(VIN), .ZN(n2120)
         );
  OAI22_X1 U2622 ( .A1(n3435), .A2(n2223), .B1(reg3_reg[1]), .B2(VIN), .ZN(
        n2119) );
  OAI22_X1 U2616 ( .A1(n3435), .A2(n2222), .B1(reg4_reg[1]), .B2(VIN), .ZN(
        n2117) );
  AOI22_X1 U2351 ( .A1(VIN), .A2(n2860), .B1(n2859), .B2(n3435), .ZN(n2414) );
  AOI22_X1 U2349 ( .A1(VIN), .A2(n2859), .B1(n2879), .B2(n3435), .ZN(n2413) );
  AOI22_X1 U2347 ( .A1(VIN), .A2(n2879), .B1(n2804), .B2(n3435), .ZN(n2412) );
  NAND2_X1 U2312 ( .A1(VIN), .A2(ff[3]), .ZN(n2008) );
  OAI21_X1 U2311 ( .B1(VIN), .B2(n2138), .A(n2008), .ZN(n2394) );
  OAI21_X1 U2636 ( .B1(VIN), .B2(n2839), .A(n2125), .ZN(n2560) );
  OAI21_X1 U2642 ( .B1(VIN), .B2(n2837), .A(n2125), .ZN(n2563) );
  OAI21_X1 U2640 ( .B1(VIN), .B2(n2868), .A(n2125), .ZN(n2562) );
  NAND2_X1 U2630 ( .A1(VIN), .A2(w[1]), .ZN(n2122) );
  OAI21_X1 U2627 ( .B1(VIN), .B2(p11_minus_A_shifted_14_), .A(n2122), .ZN(
        n2556) );
  NAND2_X1 U2599 ( .A1(VIN), .A2(w[3]), .ZN(n2113) );
  OAI21_X1 U2598 ( .B1(VIN), .B2(p11_minus_A_shifted_16_), .A(n2113), .ZN(
        n2540) );
  NAND2_X1 U2648 ( .A1(VIN), .A2(w[0]), .ZN(n2127) );
  OAI21_X1 U2645 ( .B1(VIN), .B2(n2838), .A(n2127), .ZN(n2564) );
  OAI21_X1 U2647 ( .B1(VIN), .B2(n2836), .A(n2127), .ZN(n2565) );
  OAI21_X1 U2629 ( .B1(VIN), .B2(n2864), .A(n2122), .ZN(n2557) );
  NAND2_X1 U2612 ( .A1(VIN), .A2(w[2]), .ZN(n2116) );
  OAI21_X1 U2611 ( .B1(VIN), .B2(n2820), .A(n2116), .ZN(n2548) );
  NAND2_X1 U2318 ( .A1(VIN), .A2(ff[0]), .ZN(n2011) );
  OAI21_X1 U2317 ( .B1(VIN), .B2(n2141), .A(n2011), .ZN(n2397) );
  NAND2_X1 U2314 ( .A1(VIN), .A2(ff[2]), .ZN(n2009) );
  OAI21_X1 U2313 ( .B1(VIN), .B2(n2139), .A(n2009), .ZN(n2395) );
  NAND2_X1 U2316 ( .A1(VIN), .A2(ff[1]), .ZN(n2010) );
  OAI21_X1 U2315 ( .B1(VIN), .B2(n2140), .A(n2010), .ZN(n2396) );
  NAND2_X1 U2643 ( .A1(reg2[0]), .A2(VIN), .ZN(n2125) );
  MUX2_X1 U2584 ( .A(reg2_reg[4]), .B(reg2[4]), .S(VIN), .Z(n2531) );
  MUX2_X1 U2576 ( .A(reg4_reg[4]), .B(n2216), .S(VIN), .Z(n2526) );
  MUX2_X1 U2581 ( .A(reg3_reg[4]), .B(n2217), .S(VIN), .Z(n2529) );
  NAND2_X1 U1392 ( .A1(reg1_reg[13]), .A2(n1236), .ZN(n993) );
  NAND2_X1 U1444 ( .A1(reg1_reg[11]), .A2(n1274), .ZN(n1074) );
  NAND2_X1 U640 ( .A1(reg3_reg[13]), .A2(n584), .ZN(n341) );
  NAND2_X1 U692 ( .A1(reg3_reg[11]), .A2(n622), .ZN(n422) );
  NAND2_X1 U264 ( .A1(reg4_reg[13]), .A2(n258), .ZN(n14) );
  NAND2_X1 U316 ( .A1(reg4_reg[11]), .A2(n296), .ZN(n96) );
  NAND2_X1 U1016 ( .A1(reg2_reg[13]), .A2(n910), .ZN(n667) );
  NAND2_X1 U1068 ( .A1(reg2_reg[11]), .A2(n948), .ZN(n748) );
  NAND2_X1 U1765 ( .A1(n1577), .A2(n1576), .ZN(n1411) );
  NAND2_X1 U1764 ( .A1(A1[13]), .A2(n1576), .ZN(n1412) );
  NAND2_X1 U2132 ( .A1(n1917), .A2(n1916), .ZN(n1751) );
  NAND2_X1 U2131 ( .A1(A2[13]), .A2(n1916), .ZN(n1752) );
  NAND2_X1 U1396 ( .A1(reg1_reg[11]), .A2(reg1_reg[12]), .ZN(n994) );
  NAND2_X1 U1492 ( .A1(reg1_reg[9]), .A2(n1306), .ZN(n1089) );
  NAND2_X1 U644 ( .A1(reg3_reg[11]), .A2(reg3_reg[12]), .ZN(n342) );
  NAND2_X1 U740 ( .A1(reg3_reg[9]), .A2(n654), .ZN(n437) );
  NAND2_X1 U268 ( .A1(reg4_reg[11]), .A2(reg4_reg[12]), .ZN(n15) );
  NAND2_X1 U364 ( .A1(reg4_reg[9]), .A2(n328), .ZN(n111) );
  NAND2_X1 U1020 ( .A1(reg2_reg[11]), .A2(reg2_reg[12]), .ZN(n668) );
  NAND2_X1 U1116 ( .A1(reg2_reg[9]), .A2(n980), .ZN(n763) );
  NAND2_X1 U1461 ( .A1(reg1_reg[9]), .A2(reg1_reg[10]), .ZN(n1075) );
  NAND2_X1 U709 ( .A1(reg3_reg[9]), .A2(reg3_reg[10]), .ZN(n423) );
  NAND2_X1 U333 ( .A1(reg4_reg[9]), .A2(reg4_reg[10]), .ZN(n97) );
  NAND2_X1 U1085 ( .A1(reg2_reg[9]), .A2(reg2_reg[10]), .ZN(n749) );
  NAND2_X1 U1499 ( .A1(reg1_reg[8]), .A2(p6_Partial_products_sum_add_23_B_0_), 
        .ZN(n1090) );
  NAND2_X1 U747 ( .A1(reg3_reg[8]), .A2(p8_Partial_products_sum_add_23_B_0_), 
        .ZN(n438) );
  NAND2_X1 U371 ( .A1(reg4_reg[8]), .A2(p9_Partial_products_sum_add_23_B_0_), 
        .ZN(n112) );
  NAND2_X1 U1123 ( .A1(reg2_reg[8]), .A2(p7_Partial_products_sum_add_23_B_0_), 
        .ZN(n764) );
  NAND2_X1 U1763 ( .A1(A1[13]), .A2(n1575), .ZN(n1319) );
  NAND2_X1 U2130 ( .A1(A2[13]), .A2(n1915), .ZN(n1658) );
  NAND2_X1 U2182 ( .A1(A2[11]), .A2(n1953), .ZN(n1743) );
  NAND2_X1 U1815 ( .A1(A1[11]), .A2(n1613), .ZN(n1403) );
  INV_X1 U1769 ( .A(A1[13]), .ZN(n1577) );
  INV_X1 U1813 ( .A(A1[11]), .ZN(n1578) );
  INV_X1 U1788 ( .A(A1[12]), .ZN(n1579) );
  NAND2_X1 U1768 ( .A1(A1[11]), .A2(A1[12]), .ZN(n1321) );
  INV_X1 U1767 ( .A(n1321), .ZN(n1326) );
  INV_X1 U1737 ( .A(n1411), .ZN(n1323) );
  INV_X1 U1736 ( .A(n1412), .ZN(n1324) );
  INV_X1 U1535 ( .A(p11_C[72]), .ZN(p11_S[72]) );
  INV_X1 U1863 ( .A(A1[9]), .ZN(n1394) );
  INV_X1 U1582 ( .A(n1416), .ZN(n1414) );
  INV_X1 U1762 ( .A(n1319), .ZN(n1409) );
  INV_X1 U1593 ( .A(n1333), .ZN(n1336) );
  INV_X1 U1602 ( .A(p11_muxs_out_3__20_), .ZN(n1433) );
  INV_X1 U1592 ( .A(n1426), .ZN(n1425) );
  INV_X1 U1540 ( .A(n1335), .ZN(n1334) );
  INV_X1 U1612 ( .A(n1445), .ZN(n1444) );
  INV_X1 U1609 ( .A(p11_muxs_out_3__19_), .ZN(n1345) );
  INV_X1 U1635 ( .A(p11_muxs_out_2__18_), .ZN(n1461) );
  INV_X1 U1607 ( .A(n1343), .ZN(n1344) );
  INV_X1 U1642 ( .A(p11_muxs_out_3__17_), .ZN(n1468) );
  INV_X1 U1670 ( .A(p11_muxs_out_1__16_), .ZN(n1490) );
  INV_X1 U1677 ( .A(p11_muxs_out_1__15_), .ZN(n1498) );
  INV_X1 U1657 ( .A(n1483), .ZN(n1482) );
  NOR2_X1 U1894 ( .A1(A1[1]), .A2(n1657), .ZN(n1549) );
  INV_X1 U1892 ( .A(n1590), .ZN(n1569) );
  INV_X1 U1696 ( .A(n1518), .ZN(n1515) );
  INV_X1 U1694 ( .A(n1514), .ZN(n1362) );
  INV_X1 U1884 ( .A(n1567), .ZN(n1608) );
  INV_X1 U1717 ( .A(n1538), .ZN(n1536) );
  INV_X1 U1804 ( .A(p11_muxs_out_2__11_), .ZN(n1595) );
  INV_X1 U1805 ( .A(n1596), .ZN(n1609) );
  INV_X1 U1828 ( .A(p11_muxs_out_3__10_), .ZN(n1615) );
  INV_X1 U1850 ( .A(p11_muxs_out_1__9_), .ZN(n1623) );
  INV_X1 U1851 ( .A(p11_muxs_out_2__9_), .ZN(n1624) );
  INV_X1 U1844 ( .A(n1635), .ZN(n1634) );
  INV_X1 U1837 ( .A(n1629), .ZN(n1628) );
  INV_X1 U1877 ( .A(p11_muxs_out_1__6_), .ZN(n1650) );
  INV_X1 U1873 ( .A(p11_muxs_out_3__7_), .ZN(n1399) );
  INV_X1 U1572 ( .A(n1398), .ZN(n1397) );
  INV_X1 U1896 ( .A(p11_muxs_out_3__6_), .ZN(n1654) );
  INV_X1 U2136 ( .A(A2[13]), .ZN(n1917) );
  INV_X1 U2180 ( .A(A2[11]), .ZN(n1918) );
  INV_X1 U2155 ( .A(A2[12]), .ZN(n1919) );
  NAND2_X1 U2135 ( .A1(A2[11]), .A2(A2[12]), .ZN(n1660) );
  INV_X1 U2134 ( .A(n1660), .ZN(n1665) );
  INV_X1 U2104 ( .A(n1751), .ZN(n1662) );
  INV_X1 U2103 ( .A(n1752), .ZN(n1663) );
  INV_X1 U1902 ( .A(p10_C[72]), .ZN(p10_S[72]) );
  NAND2_X1 U2227 ( .A1(A2[9]), .A2(n1985), .ZN(n1760) );
  INV_X1 U2230 ( .A(A2[9]), .ZN(n1734) );
  INV_X1 U1949 ( .A(n1756), .ZN(n1754) );
  INV_X1 U2129 ( .A(n1658), .ZN(n1749) );
  INV_X1 U1960 ( .A(n1673), .ZN(n1676) );
  INV_X1 U1969 ( .A(p10_muxs_out_3__20_), .ZN(n1773) );
  INV_X1 U1959 ( .A(n1766), .ZN(n1765) );
  INV_X1 U1907 ( .A(n1675), .ZN(n1674) );
  INV_X1 U1979 ( .A(n1785), .ZN(n1784) );
  INV_X1 U1976 ( .A(p10_muxs_out_3__19_), .ZN(n1685) );
  INV_X1 U2002 ( .A(p10_muxs_out_2__18_), .ZN(n1801) );
  INV_X1 U1974 ( .A(n1683), .ZN(n1684) );
  INV_X1 U2009 ( .A(p10_muxs_out_3__17_), .ZN(n1808) );
  INV_X1 U2037 ( .A(p10_muxs_out_1__16_), .ZN(n1830) );
  INV_X1 U2044 ( .A(p10_muxs_out_1__15_), .ZN(n1838) );
  INV_X1 U2024 ( .A(n1823), .ZN(n1822) );
  INV_X1 U2262 ( .A(A2[0]), .ZN(n1997) );
  NOR2_X1 U2261 ( .A1(A2[1]), .A2(n1997), .ZN(n1889) );
  INV_X1 U2259 ( .A(n1930), .ZN(n1909) );
  INV_X1 U2063 ( .A(n1858), .ZN(n1855) );
  INV_X1 U2061 ( .A(n1854), .ZN(n1702) );
  INV_X1 U2251 ( .A(n1907), .ZN(n1948) );
  INV_X1 U2084 ( .A(n1878), .ZN(n1876) );
  INV_X1 U2171 ( .A(p10_muxs_out_2__11_), .ZN(n1935) );
  INV_X1 U2172 ( .A(n1936), .ZN(n1949) );
  INV_X1 U2194 ( .A(p10_muxs_out_2__10_), .ZN(n1954) );
  INV_X1 U2195 ( .A(p10_muxs_out_3__10_), .ZN(n1955) );
  INV_X1 U2217 ( .A(p10_muxs_out_1__9_), .ZN(n1963) );
  INV_X1 U2218 ( .A(p10_muxs_out_2__9_), .ZN(n1964) );
  INV_X1 U2228 ( .A(n1770), .ZN(n1973) );
  INV_X1 U2211 ( .A(n1975), .ZN(n1974) );
  INV_X1 U2204 ( .A(n1969), .ZN(n1968) );
  INV_X1 U2244 ( .A(p10_muxs_out_1__6_), .ZN(n1990) );
  INV_X1 U2240 ( .A(p10_muxs_out_3__7_), .ZN(n1739) );
  INV_X1 U1939 ( .A(n1738), .ZN(n1737) );
  INV_X1 U2263 ( .A(p10_muxs_out_3__6_), .ZN(n1994) );
  INV_X1 U1407 ( .A(B0[12]), .ZN(p6_minus_A_shifted_25_) );
  INV_X1 U1155 ( .A(p6_final_product2_26_), .ZN(p6_final_product2_25_) );
  INV_X1 U1159 ( .A(p6_C[72]), .ZN(p6_S[72]) );
  INV_X1 U1206 ( .A(n1086), .ZN(n1084) );
  INV_X1 U1249 ( .A(n994), .ZN(n998) );
  INV_X1 U1250 ( .A(n993), .ZN(n1079) );
  INV_X1 U1368 ( .A(n996), .ZN(n1081) );
  INV_X1 U1369 ( .A(n997), .ZN(n1082) );
  INV_X1 U1217 ( .A(n1005), .ZN(n1008) );
  INV_X1 U1226 ( .A(p6_muxs_out_3__20_), .ZN(n1102) );
  INV_X1 U1216 ( .A(n1095), .ZN(n1094) );
  INV_X1 U1164 ( .A(n1007), .ZN(n1006) );
  INV_X1 U1236 ( .A(n1113), .ZN(n1112) );
  INV_X1 U1233 ( .A(p6_muxs_out_3__19_), .ZN(n1017) );
  INV_X1 U1262 ( .A(p6_muxs_out_2__18_), .ZN(n1127) );
  INV_X1 U1231 ( .A(n1015), .ZN(n1016) );
  INV_X1 U1269 ( .A(p6_muxs_out_3__17_), .ZN(n1134) );
  INV_X1 U1297 ( .A(p6_muxs_out_1__16_), .ZN(n1154) );
  INV_X1 U1304 ( .A(p6_muxs_out_1__15_), .ZN(n1162) );
  INV_X1 U1284 ( .A(n1148), .ZN(n1147) );
  INV_X1 U1464 ( .A(B0[2]), .ZN(p6_minus_A_shifted_15_) );
  INV_X1 U1526 ( .A(n1246), .ZN(n1230) );
  INV_X1 U1476 ( .A(B0[1]), .ZN(p6_minus_A_shifted_14_) );
  INV_X1 U1517 ( .A(n1212), .ZN(n1247) );
  INV_X1 U1323 ( .A(n1181), .ZN(n1178) );
  INV_X1 U1321 ( .A(n1177), .ZN(n1034) );
  INV_X1 U1495 ( .A(B0[0]), .ZN(p6_minus_A_shifted_13_) );
  INV_X1 U1518 ( .A(n1228), .ZN(n1269) );
  INV_X1 U1345 ( .A(n1201), .ZN(n1198) );
  INV_X1 U1343 ( .A(n1197), .ZN(n1038) );
  INV_X1 U1433 ( .A(p6_muxs_out_2__11_), .ZN(n1255) );
  INV_X1 U1434 ( .A(n1256), .ZN(n1270) );
  INV_X1 U1456 ( .A(p6_muxs_out_2__10_), .ZN(n1275) );
  INV_X1 U1457 ( .A(p6_muxs_out_3__10_), .ZN(n1276) );
  INV_X1 U1483 ( .A(p6_muxs_out_2__9_), .ZN(n1285) );
  INV_X1 U1482 ( .A(p6_muxs_out_1__9_), .ZN(n1284) );
  INV_X1 U1496 ( .A(n1098), .ZN(n1293) );
  INV_X1 U1493 ( .A(n1099), .ZN(n1294) );
  INV_X1 U1474 ( .A(n1296), .ZN(n1295) );
  INV_X1 U1467 ( .A(n1290), .ZN(n1289) );
  INV_X1 U1510 ( .A(p6_muxs_out_1__6_), .ZN(n1311) );
  INV_X1 U1530 ( .A(p6_muxs_out_3__6_), .ZN(n1315) );
  INV_X1 U1196 ( .A(n1070), .ZN(n1069) );
  INV_X1 U1506 ( .A(p6_muxs_out_3__7_), .ZN(n1071) );
  INV_X1 U497 ( .A(n342), .ZN(n346) );
  INV_X1 U655 ( .A(B2[12]), .ZN(p8_minus_A_shifted_25_) );
  INV_X1 U403 ( .A(p8_final_product2_26_), .ZN(p8_final_product2_25_) );
  INV_X1 U407 ( .A(p8_C[72]), .ZN(p8_S[72]) );
  INV_X1 U454 ( .A(n434), .ZN(n432) );
  INV_X1 U498 ( .A(n341), .ZN(n427) );
  INV_X1 U616 ( .A(n344), .ZN(n429) );
  INV_X1 U617 ( .A(n345), .ZN(n430) );
  INV_X1 U465 ( .A(n353), .ZN(n356) );
  INV_X1 U474 ( .A(p8_muxs_out_3__20_), .ZN(n450) );
  INV_X1 U464 ( .A(n443), .ZN(n442) );
  INV_X1 U412 ( .A(n355), .ZN(n354) );
  INV_X1 U484 ( .A(n461), .ZN(n460) );
  INV_X1 U481 ( .A(p8_muxs_out_3__19_), .ZN(n365) );
  INV_X1 U510 ( .A(p8_muxs_out_2__18_), .ZN(n475) );
  INV_X1 U479 ( .A(n363), .ZN(n364) );
  INV_X1 U517 ( .A(p8_muxs_out_3__17_), .ZN(n482) );
  INV_X1 U545 ( .A(p8_muxs_out_1__16_), .ZN(n502) );
  INV_X1 U552 ( .A(p8_muxs_out_1__15_), .ZN(n510) );
  INV_X1 U532 ( .A(n496), .ZN(n495) );
  INV_X1 U686 ( .A(B2[3]), .ZN(p8_minus_A_shifted_16_) );
  INV_X1 U712 ( .A(B2[2]), .ZN(p8_minus_A_shifted_15_) );
  INV_X1 U774 ( .A(n594), .ZN(n578) );
  INV_X1 U765 ( .A(n560), .ZN(n595) );
  INV_X1 U571 ( .A(n529), .ZN(n526) );
  INV_X1 U569 ( .A(n525), .ZN(n382) );
  INV_X1 U743 ( .A(B2[0]), .ZN(p8_minus_A_shifted_13_) );
  INV_X1 U766 ( .A(n576), .ZN(n617) );
  INV_X1 U593 ( .A(n549), .ZN(n546) );
  INV_X1 U591 ( .A(n545), .ZN(n386) );
  INV_X1 U681 ( .A(p8_muxs_out_2__11_), .ZN(n603) );
  INV_X1 U682 ( .A(n604), .ZN(n618) );
  INV_X1 U704 ( .A(p8_muxs_out_2__10_), .ZN(n623) );
  INV_X1 U705 ( .A(p8_muxs_out_3__10_), .ZN(n624) );
  INV_X1 U730 ( .A(p8_muxs_out_1__9_), .ZN(n632) );
  INV_X1 U731 ( .A(p8_muxs_out_2__9_), .ZN(n633) );
  INV_X1 U744 ( .A(n446), .ZN(n641) );
  INV_X1 U741 ( .A(n447), .ZN(n642) );
  INV_X1 U722 ( .A(n644), .ZN(n643) );
  INV_X1 U715 ( .A(n638), .ZN(n637) );
  INV_X1 U758 ( .A(p8_muxs_out_1__6_), .ZN(n659) );
  INV_X1 U441 ( .A(n413), .ZN(n412) );
  INV_X1 U754 ( .A(p8_muxs_out_3__7_), .ZN(n419) );
  INV_X1 U444 ( .A(n418), .ZN(n417) );
  INV_X1 U778 ( .A(p8_muxs_out_3__6_), .ZN(n663) );
  INV_X1 U121 ( .A(n15), .ZN(n20) );
  INV_X1 U279 ( .A(B3[12]), .ZN(p9_minus_A_shifted_25_) );
  INV_X1 U3 ( .A(p9_final_product2_26_), .ZN(p9_final_product2_25_) );
  INV_X1 U25 ( .A(p9_C[72]), .ZN(p9_S[72]) );
  INV_X1 U78 ( .A(n108), .ZN(n106) );
  INV_X1 U122 ( .A(n14), .ZN(n101) );
  INV_X1 U240 ( .A(n17), .ZN(n103) );
  INV_X1 U241 ( .A(n18), .ZN(n104) );
  INV_X1 U89 ( .A(n27), .ZN(n30) );
  INV_X1 U98 ( .A(p9_muxs_out_3__20_), .ZN(n124) );
  INV_X1 U88 ( .A(n117), .ZN(n116) );
  INV_X1 U30 ( .A(n29), .ZN(n28) );
  INV_X1 U108 ( .A(n135), .ZN(n134) );
  INV_X1 U105 ( .A(p9_muxs_out_3__19_), .ZN(n39) );
  INV_X1 U134 ( .A(p9_muxs_out_2__18_), .ZN(n149) );
  INV_X1 U103 ( .A(n37), .ZN(n38) );
  INV_X1 U141 ( .A(p9_muxs_out_3__17_), .ZN(n156) );
  INV_X1 U169 ( .A(p9_muxs_out_1__16_), .ZN(n176) );
  INV_X1 U176 ( .A(p9_muxs_out_1__15_), .ZN(n184) );
  INV_X1 U156 ( .A(n170), .ZN(n169) );
  INV_X1 U310 ( .A(B3[3]), .ZN(p9_minus_A_shifted_16_) );
  INV_X1 U336 ( .A(B3[2]), .ZN(p9_minus_A_shifted_15_) );
  INV_X1 U398 ( .A(n268), .ZN(n252) );
  INV_X1 U389 ( .A(n234), .ZN(n269) );
  INV_X1 U195 ( .A(n203), .ZN(n200) );
  INV_X1 U193 ( .A(n199), .ZN(n56) );
  INV_X1 U367 ( .A(B3[0]), .ZN(p9_minus_A_shifted_13_) );
  INV_X1 U390 ( .A(n250), .ZN(n291) );
  INV_X1 U217 ( .A(n223), .ZN(n220) );
  INV_X1 U215 ( .A(n219), .ZN(n60) );
  INV_X1 U305 ( .A(p9_muxs_out_2__11_), .ZN(n277) );
  INV_X1 U306 ( .A(n278), .ZN(n292) );
  INV_X1 U328 ( .A(p9_muxs_out_2__10_), .ZN(n297) );
  INV_X1 U329 ( .A(p9_muxs_out_3__10_), .ZN(n298) );
  INV_X1 U354 ( .A(p9_muxs_out_1__9_), .ZN(n306) );
  INV_X1 U355 ( .A(p9_muxs_out_2__9_), .ZN(n307) );
  INV_X1 U368 ( .A(n120), .ZN(n315) );
  INV_X1 U365 ( .A(n121), .ZN(n316) );
  INV_X1 U346 ( .A(n318), .ZN(n317) );
  INV_X1 U339 ( .A(n312), .ZN(n311) );
  INV_X1 U382 ( .A(p9_muxs_out_1__6_), .ZN(n333) );
  INV_X1 U65 ( .A(n87), .ZN(n86) );
  INV_X1 U378 ( .A(p9_muxs_out_3__7_), .ZN(n93) );
  INV_X1 U68 ( .A(n92), .ZN(n91) );
  INV_X1 U402 ( .A(p9_muxs_out_3__6_), .ZN(n337) );
  INV_X1 U873 ( .A(n668), .ZN(n672) );
  INV_X1 U1031 ( .A(B1[12]), .ZN(p7_minus_A_shifted_25_) );
  INV_X1 U779 ( .A(p7_final_product2_26_), .ZN(p7_final_product2_25_) );
  INV_X1 U783 ( .A(p7_C[72]), .ZN(p7_S[72]) );
  INV_X1 U830 ( .A(n760), .ZN(n758) );
  INV_X1 U874 ( .A(n667), .ZN(n753) );
  INV_X1 U992 ( .A(n670), .ZN(n755) );
  INV_X1 U993 ( .A(n671), .ZN(n756) );
  INV_X1 U841 ( .A(n679), .ZN(n682) );
  INV_X1 U850 ( .A(p7_muxs_out_3__20_), .ZN(n776) );
  INV_X1 U840 ( .A(n769), .ZN(n768) );
  INV_X1 U788 ( .A(n681), .ZN(n680) );
  INV_X1 U860 ( .A(n787), .ZN(n786) );
  INV_X1 U857 ( .A(p7_muxs_out_3__19_), .ZN(n691) );
  INV_X1 U886 ( .A(p7_muxs_out_2__18_), .ZN(n801) );
  INV_X1 U855 ( .A(n689), .ZN(n690) );
  INV_X1 U893 ( .A(p7_muxs_out_3__17_), .ZN(n808) );
  INV_X1 U921 ( .A(p7_muxs_out_1__16_), .ZN(n828) );
  INV_X1 U928 ( .A(p7_muxs_out_1__15_), .ZN(n836) );
  INV_X1 U908 ( .A(n822), .ZN(n821) );
  INV_X1 U1062 ( .A(B1[3]), .ZN(p7_minus_A_shifted_16_) );
  INV_X1 U1088 ( .A(B1[2]), .ZN(p7_minus_A_shifted_15_) );
  INV_X1 U1150 ( .A(n920), .ZN(n904) );
  INV_X1 U1141 ( .A(n886), .ZN(n921) );
  INV_X1 U947 ( .A(n855), .ZN(n852) );
  INV_X1 U945 ( .A(n851), .ZN(n708) );
  INV_X1 U1119 ( .A(B1[0]), .ZN(p7_minus_A_shifted_13_) );
  INV_X1 U1142 ( .A(n902), .ZN(n943) );
  INV_X1 U969 ( .A(n875), .ZN(n872) );
  INV_X1 U967 ( .A(n871), .ZN(n712) );
  INV_X1 U1057 ( .A(p7_muxs_out_2__11_), .ZN(n929) );
  INV_X1 U1058 ( .A(n930), .ZN(n944) );
  INV_X1 U1080 ( .A(p7_muxs_out_2__10_), .ZN(n949) );
  INV_X1 U1081 ( .A(p7_muxs_out_3__10_), .ZN(n950) );
  INV_X1 U1106 ( .A(p7_muxs_out_1__9_), .ZN(n958) );
  INV_X1 U1107 ( .A(p7_muxs_out_2__9_), .ZN(n959) );
  INV_X1 U1120 ( .A(n772), .ZN(n967) );
  INV_X1 U1117 ( .A(n773), .ZN(n968) );
  INV_X1 U1098 ( .A(n970), .ZN(n969) );
  INV_X1 U1091 ( .A(n964), .ZN(n963) );
  INV_X1 U1134 ( .A(p7_muxs_out_1__6_), .ZN(n985) );
  INV_X1 U817 ( .A(n739), .ZN(n738) );
  INV_X1 U1130 ( .A(p7_muxs_out_3__7_), .ZN(n745) );
  INV_X1 U820 ( .A(n744), .ZN(n743) );
  INV_X1 U1154 ( .A(p7_muxs_out_3__6_), .ZN(n989) );
  INV_X1 U2617 ( .A(n2118), .ZN(n2551) );
  INV_X1 U2623 ( .A(n2120), .ZN(n2554) );
  INV_X1 U2621 ( .A(n2119), .ZN(n2553) );
  INV_X1 U2615 ( .A(n2117), .ZN(n2550) );
  HA_X1 s8_add_23_DP_OP_277_3998_2_U48 ( .A(mul3_reg[0]), .B(mul2_reg[0]), 
        .CO(s8_add_23_DP_OP_277_3998_2_n90), .S(s8_add_23_DP_OP_277_3998_2_n91) );
  HA_X1 s8_add_23_DP_OP_277_3998_2_U47 ( .A(mul4_reg[1]), .B(mul2_reg[1]), 
        .CO(s8_add_23_DP_OP_277_3998_2_n88), .S(s8_add_23_DP_OP_277_3998_2_n89) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U46 ( .A(mul1_reg[1]), .B(mul3_reg[1]), 
        .CI(s8_add_23_DP_OP_277_3998_2_n90), .CO(
        s8_add_23_DP_OP_277_3998_2_n86), .S(s8_add_23_DP_OP_277_3998_2_n87) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U45 ( .A(mul4_reg[2]), .B(mul2_reg[2]), 
        .CI(mul1_reg[2]), .CO(s8_add_23_DP_OP_277_3998_2_n84), .S(
        s8_add_23_DP_OP_277_3998_2_n85) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U44 ( .A(s8_add_23_DP_OP_277_3998_2_n88), 
        .B(mul3_reg[2]), .CI(s8_add_23_DP_OP_277_3998_2_n86), .CO(
        s8_add_23_DP_OP_277_3998_2_n82), .S(s8_add_23_DP_OP_277_3998_2_n83) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U43 ( .A(mul4_reg[3]), .B(mul2_reg[3]), 
        .CI(mul1_reg[3]), .CO(s8_add_23_DP_OP_277_3998_2_n80), .S(
        s8_add_23_DP_OP_277_3998_2_n81) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U42 ( .A(s8_add_23_DP_OP_277_3998_2_n84), 
        .B(mul3_reg[3]), .CI(s8_add_23_DP_OP_277_3998_2_n81), .CO(
        s8_add_23_DP_OP_277_3998_2_n78), .S(s8_add_23_DP_OP_277_3998_2_n79) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U41 ( .A(mul4_reg[4]), .B(mul2_reg[4]), 
        .CI(mul1_reg[4]), .CO(s8_add_23_DP_OP_277_3998_2_n76), .S(
        s8_add_23_DP_OP_277_3998_2_n77) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U40 ( .A(s8_add_23_DP_OP_277_3998_2_n80), 
        .B(mul3_reg[4]), .CI(s8_add_23_DP_OP_277_3998_2_n77), .CO(
        s8_add_23_DP_OP_277_3998_2_n74), .S(s8_add_23_DP_OP_277_3998_2_n75) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U39 ( .A(mul4_reg[5]), .B(mul2_reg[5]), 
        .CI(mul1_reg[5]), .CO(s8_add_23_DP_OP_277_3998_2_n72), .S(
        s8_add_23_DP_OP_277_3998_2_n73) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U38 ( .A(s8_add_23_DP_OP_277_3998_2_n76), 
        .B(mul3_reg[5]), .CI(s8_add_23_DP_OP_277_3998_2_n73), .CO(
        s8_add_23_DP_OP_277_3998_2_n70), .S(s8_add_23_DP_OP_277_3998_2_n71) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U37 ( .A(mul4_reg[6]), .B(mul2_reg[6]), 
        .CI(mul1_reg[6]), .CO(s8_add_23_DP_OP_277_3998_2_n68), .S(
        s8_add_23_DP_OP_277_3998_2_n69) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U36 ( .A(s8_add_23_DP_OP_277_3998_2_n72), 
        .B(mul3_reg[6]), .CI(s8_add_23_DP_OP_277_3998_2_n69), .CO(
        s8_add_23_DP_OP_277_3998_2_n66), .S(s8_add_23_DP_OP_277_3998_2_n67) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U35 ( .A(mul4_reg[7]), .B(mul2_reg[7]), 
        .CI(mul1_reg[7]), .CO(s8_add_23_DP_OP_277_3998_2_n64), .S(
        s8_add_23_DP_OP_277_3998_2_n65) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U34 ( .A(s8_add_23_DP_OP_277_3998_2_n68), 
        .B(mul3_reg[7]), .CI(s8_add_23_DP_OP_277_3998_2_n65), .CO(
        s8_add_23_DP_OP_277_3998_2_n62), .S(s8_add_23_DP_OP_277_3998_2_n63) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U33 ( .A(mul4_reg[8]), .B(mul2_reg[8]), 
        .CI(mul1_reg[8]), .CO(s8_add_23_DP_OP_277_3998_2_n60), .S(
        s8_add_23_DP_OP_277_3998_2_n61) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U32 ( .A(s8_add_23_DP_OP_277_3998_2_n64), 
        .B(mul3_reg[8]), .CI(s8_add_23_DP_OP_277_3998_2_n61), .CO(
        s8_add_23_DP_OP_277_3998_2_n58), .S(s8_add_23_DP_OP_277_3998_2_n59) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U31 ( .A(mul4_reg[9]), .B(mul2_reg[9]), 
        .CI(mul1_reg[9]), .CO(s8_add_23_DP_OP_277_3998_2_n56), .S(
        s8_add_23_DP_OP_277_3998_2_n57) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U30 ( .A(s8_add_23_DP_OP_277_3998_2_n60), 
        .B(mul3_reg[9]), .CI(s8_add_23_DP_OP_277_3998_2_n57), .CO(
        s8_add_23_DP_OP_277_3998_2_n54), .S(s8_add_23_DP_OP_277_3998_2_n55) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U29 ( .A(mul4_reg[10]), .B(mul2_reg[10]), 
        .CI(mul1_reg[10]), .CO(s8_add_23_DP_OP_277_3998_2_n52), .S(
        s8_add_23_DP_OP_277_3998_2_n53) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U28 ( .A(s8_add_23_DP_OP_277_3998_2_n56), 
        .B(mul3_reg[10]), .CI(s8_add_23_DP_OP_277_3998_2_n53), .CO(
        s8_add_23_DP_OP_277_3998_2_n50), .S(s8_add_23_DP_OP_277_3998_2_n51) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U27 ( .A(mul4_reg[11]), .B(mul2_reg[11]), 
        .CI(mul1_reg[11]), .CO(s8_add_23_DP_OP_277_3998_2_n48), .S(
        s8_add_23_DP_OP_277_3998_2_n49) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U26 ( .A(s8_add_23_DP_OP_277_3998_2_n52), 
        .B(mul3_reg[11]), .CI(s8_add_23_DP_OP_277_3998_2_n49), .CO(
        s8_add_23_DP_OP_277_3998_2_n46), .S(s8_add_23_DP_OP_277_3998_2_n47) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U25 ( .A(mul4_reg[12]), .B(mul2_reg[12]), 
        .CI(mul1_reg[12]), .CO(s8_add_23_DP_OP_277_3998_2_n44), .S(
        s8_add_23_DP_OP_277_3998_2_n45) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U24 ( .A(s8_add_23_DP_OP_277_3998_2_n48), 
        .B(mul3_reg[12]), .CI(s8_add_23_DP_OP_277_3998_2_n45), .CO(
        s8_add_23_DP_OP_277_3998_2_n42), .S(s8_add_23_DP_OP_277_3998_2_n43) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U23 ( .A(mul4_reg[0]), .B(mul1_reg[0]), 
        .CI(s8_add_23_DP_OP_277_3998_2_n91), .CO(
        s8_add_23_DP_OP_277_3998_2_n39), .S(ff[0]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U20 ( .A(s8_add_23_DP_OP_277_3998_2_n39), 
        .B(s8_add_23_DP_OP_277_3998_2_n89), .CI(s8_add_23_DP_OP_277_3998_2_n87), .CO(s8_add_23_DP_OP_277_3998_2_n38), .S(ff[1]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U19 ( .A(s8_add_23_DP_OP_277_3998_2_n83), 
        .B(s8_add_23_DP_OP_277_3998_2_n85), .CI(s8_add_23_DP_OP_277_3998_2_n38), .CO(s8_add_23_DP_OP_277_3998_2_n37), .S(ff[2]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U18 ( .A(s8_add_23_DP_OP_277_3998_2_n79), 
        .B(s8_add_23_DP_OP_277_3998_2_n82), .CI(s8_add_23_DP_OP_277_3998_2_n37), .CO(s8_add_23_DP_OP_277_3998_2_n36), .S(ff[3]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U17 ( .A(s8_add_23_DP_OP_277_3998_2_n75), 
        .B(s8_add_23_DP_OP_277_3998_2_n78), .CI(s8_add_23_DP_OP_277_3998_2_n36), .CO(s8_add_23_DP_OP_277_3998_2_n35), .S(ff[4]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U16 ( .A(s8_add_23_DP_OP_277_3998_2_n71), 
        .B(s8_add_23_DP_OP_277_3998_2_n74), .CI(s8_add_23_DP_OP_277_3998_2_n35), .CO(s8_add_23_DP_OP_277_3998_2_n34), .S(ff[5]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U15 ( .A(s8_add_23_DP_OP_277_3998_2_n67), 
        .B(s8_add_23_DP_OP_277_3998_2_n70), .CI(s8_add_23_DP_OP_277_3998_2_n34), .CO(s8_add_23_DP_OP_277_3998_2_n33), .S(ff[6]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U14 ( .A(s8_add_23_DP_OP_277_3998_2_n63), 
        .B(s8_add_23_DP_OP_277_3998_2_n66), .CI(s8_add_23_DP_OP_277_3998_2_n33), .CO(s8_add_23_DP_OP_277_3998_2_n32), .S(ff[7]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U13 ( .A(s8_add_23_DP_OP_277_3998_2_n59), 
        .B(s8_add_23_DP_OP_277_3998_2_n62), .CI(s8_add_23_DP_OP_277_3998_2_n32), .CO(s8_add_23_DP_OP_277_3998_2_n31), .S(ff[8]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U10 ( .A(s8_add_23_DP_OP_277_3998_2_n55), 
        .B(s8_add_23_DP_OP_277_3998_2_n58), .CI(s8_add_23_DP_OP_277_3998_2_n31), .CO(s8_add_23_DP_OP_277_3998_2_n30), .S(ff[9]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U9 ( .A(s8_add_23_DP_OP_277_3998_2_n51), 
        .B(s8_add_23_DP_OP_277_3998_2_n54), .CI(s8_add_23_DP_OP_277_3998_2_n30), .CO(s8_add_23_DP_OP_277_3998_2_n29), .S(ff[10]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U8 ( .A(s8_add_23_DP_OP_277_3998_2_n47), 
        .B(s8_add_23_DP_OP_277_3998_2_n50), .CI(s8_add_23_DP_OP_277_3998_2_n29), .CO(s8_add_23_DP_OP_277_3998_2_n28), .S(ff[11]) );
  FA_X1 s8_add_23_DP_OP_277_3998_2_U7 ( .A(s8_add_23_DP_OP_277_3998_2_n43), 
        .B(s8_add_23_DP_OP_277_3998_2_n46), .CI(s8_add_23_DP_OP_277_3998_2_n28), .CO(s8_add_23_DP_OP_277_3998_2_n27), .S(ff[12]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U33 ( .A(n2668), .B(xin[2]), .CI(n2681), 
        .CO(s9_add_23_DP_OP_276_9387_1_n57), .S(s9_add_23_DP_OP_276_9387_1_n58) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U32 ( .A(n2667), .B(xin[3]), .CI(n2680), 
        .CO(s9_add_23_DP_OP_276_9387_1_n55), .S(s9_add_23_DP_OP_276_9387_1_n56) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U31 ( .A(n2666), .B(xin[4]), .CI(n2679), 
        .CO(s9_add_23_DP_OP_276_9387_1_n53), .S(s9_add_23_DP_OP_276_9387_1_n54) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U30 ( .A(n2665), .B(xin[5]), .CI(n2678), 
        .CO(s9_add_23_DP_OP_276_9387_1_n51), .S(s9_add_23_DP_OP_276_9387_1_n52) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U29 ( .A(n2664), .B(xin[6]), .CI(n2677), 
        .CO(s9_add_23_DP_OP_276_9387_1_n49), .S(s9_add_23_DP_OP_276_9387_1_n50) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U28 ( .A(n2663), .B(xin[7]), .CI(n2676), 
        .CO(s9_add_23_DP_OP_276_9387_1_n47), .S(s9_add_23_DP_OP_276_9387_1_n48) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U27 ( .A(n2662), .B(xin[8]), .CI(n2675), 
        .CO(s9_add_23_DP_OP_276_9387_1_n45), .S(s9_add_23_DP_OP_276_9387_1_n46) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U26 ( .A(n2661), .B(xin[9]), .CI(n2674), 
        .CO(s9_add_23_DP_OP_276_9387_1_n43), .S(s9_add_23_DP_OP_276_9387_1_n44) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U25 ( .A(n2671), .B(xin[10]), .CI(n2685), 
        .CO(s9_add_23_DP_OP_276_9387_1_n41), .S(s9_add_23_DP_OP_276_9387_1_n42) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U24 ( .A(n2670), .B(xin[11]), .CI(n2684), 
        .CO(s9_add_23_DP_OP_276_9387_1_n39), .S(s9_add_23_DP_OP_276_9387_1_n40) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U23 ( .A(n2669), .B(xin[12]), .CI(n2683), 
        .CO(s9_add_23_DP_OP_276_9387_1_n37), .S(s9_add_23_DP_OP_276_9387_1_n38) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U20 ( .A(n2660), .B(xin[0]), .CI(n2673), 
        .CO(s9_add_23_DP_OP_276_9387_1_n34), .S(w[0]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U19 ( .A(s9_add_23_DP_OP_276_9387_1_n60), 
        .B(n2672), .CI(s9_add_23_DP_OP_276_9387_1_n34), .CO(
        s9_add_23_DP_OP_276_9387_1_n33), .S(w[1]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U18 ( .A(s9_add_23_DP_OP_276_9387_1_n58), 
        .B(s9_add_23_DP_OP_276_9387_1_n59), .CI(s9_add_23_DP_OP_276_9387_1_n33), .CO(s9_add_23_DP_OP_276_9387_1_n32), .S(w[2]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U17 ( .A(s9_add_23_DP_OP_276_9387_1_n56), 
        .B(s9_add_23_DP_OP_276_9387_1_n57), .CI(s9_add_23_DP_OP_276_9387_1_n32), .CO(s9_add_23_DP_OP_276_9387_1_n31), .S(w[3]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U16 ( .A(s9_add_23_DP_OP_276_9387_1_n54), 
        .B(s9_add_23_DP_OP_276_9387_1_n55), .CI(s9_add_23_DP_OP_276_9387_1_n31), .CO(s9_add_23_DP_OP_276_9387_1_n30), .S(w[4]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U15 ( .A(s9_add_23_DP_OP_276_9387_1_n52), 
        .B(s9_add_23_DP_OP_276_9387_1_n53), .CI(s9_add_23_DP_OP_276_9387_1_n30), .CO(s9_add_23_DP_OP_276_9387_1_n29), .S(w[5]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U14 ( .A(s9_add_23_DP_OP_276_9387_1_n50), 
        .B(s9_add_23_DP_OP_276_9387_1_n51), .CI(s9_add_23_DP_OP_276_9387_1_n29), .CO(s9_add_23_DP_OP_276_9387_1_n28), .S(w[6]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U13 ( .A(s9_add_23_DP_OP_276_9387_1_n48), 
        .B(s9_add_23_DP_OP_276_9387_1_n49), .CI(s9_add_23_DP_OP_276_9387_1_n28), .CO(s9_add_23_DP_OP_276_9387_1_n27), .S(w[7]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U12 ( .A(s9_add_23_DP_OP_276_9387_1_n46), 
        .B(s9_add_23_DP_OP_276_9387_1_n47), .CI(s9_add_23_DP_OP_276_9387_1_n27), .CO(s9_add_23_DP_OP_276_9387_1_n26), .S(w[8]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U10 ( .A(s9_add_23_DP_OP_276_9387_1_n44), 
        .B(s9_add_23_DP_OP_276_9387_1_n45), .CI(s9_add_23_DP_OP_276_9387_1_n26), .CO(s9_add_23_DP_OP_276_9387_1_n25), .S(w[9]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U9 ( .A(s9_add_23_DP_OP_276_9387_1_n42), 
        .B(s9_add_23_DP_OP_276_9387_1_n43), .CI(s9_add_23_DP_OP_276_9387_1_n25), .CO(s9_add_23_DP_OP_276_9387_1_n24), .S(w[10]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U8 ( .A(s9_add_23_DP_OP_276_9387_1_n40), 
        .B(s9_add_23_DP_OP_276_9387_1_n41), .CI(s9_add_23_DP_OP_276_9387_1_n24), .CO(s9_add_23_DP_OP_276_9387_1_n23), .S(w[11]) );
  FA_X1 s9_add_23_DP_OP_276_9387_1_U7 ( .A(s9_add_23_DP_OP_276_9387_1_n38), 
        .B(s9_add_23_DP_OP_276_9387_1_n39), .CI(s9_add_23_DP_OP_276_9387_1_n23), .CO(s9_add_23_DP_OP_276_9387_1_n22), .S(w[12]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_7 ( .A(p10_S[61]), .B(p10_C[60]), 
        .CI(p10_Partial_products_sum_add_23_carry_7_), .CO(
        p10_Partial_products_sum_add_23_carry_8_), .S(temp5[0]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_8 ( .A(p10_S[62]), .B(p10_C[61]), 
        .CI(p10_Partial_products_sum_add_23_carry_8_), .CO(
        p10_Partial_products_sum_add_23_carry_9_), .S(temp5[1]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_9 ( .A(p10_S[63]), .B(p10_C[62]), 
        .CI(p10_Partial_products_sum_add_23_carry_9_), .CO(
        p10_Partial_products_sum_add_23_carry_10_), .S(temp5[2]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_10 ( .A(p10_S[64]), .B(p10_C[63]), 
        .CI(p10_Partial_products_sum_add_23_carry_10_), .CO(
        p10_Partial_products_sum_add_23_carry_11_), .S(temp5[3]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_11 ( .A(p10_S[65]), .B(p10_C[64]), 
        .CI(p10_Partial_products_sum_add_23_carry_11_), .CO(
        p10_Partial_products_sum_add_23_carry_12_), .S(temp5[4]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_12 ( .A(p10_S[66]), .B(p10_C[65]), 
        .CI(p10_Partial_products_sum_add_23_carry_12_), .CO(
        p10_Partial_products_sum_add_23_carry_13_), .S(temp5[5]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_13 ( .A(p10_S[67]), .B(p10_C[66]), 
        .CI(p10_Partial_products_sum_add_23_carry_13_), .CO(
        p10_Partial_products_sum_add_23_carry_14_), .S(temp5[6]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_14 ( .A(p10_S[68]), .B(p10_C[67]), 
        .CI(p10_Partial_products_sum_add_23_carry_14_), .CO(
        p10_Partial_products_sum_add_23_carry_15_), .S(temp5[7]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_15 ( .A(p10_S[69]), .B(p10_C[68]), 
        .CI(p10_Partial_products_sum_add_23_carry_15_), .CO(
        p10_Partial_products_sum_add_23_carry_16_), .S(temp5[8]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_16 ( .A(p10_S[70]), .B(p10_C[69]), 
        .CI(p10_Partial_products_sum_add_23_carry_16_), .CO(
        p10_Partial_products_sum_add_23_carry_17_), .S(temp5[9]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_17 ( .A(p10_S[71]), .B(p10_C[70]), 
        .CI(p10_Partial_products_sum_add_23_carry_17_), .CO(
        p10_Partial_products_sum_add_23_carry_18_), .S(temp5[10]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_18 ( .A(p10_S[72]), .B(p10_C[71]), 
        .CI(p10_Partial_products_sum_add_23_carry_18_), .CO(
        p10_Partial_products_sum_add_23_carry_19_), .S(temp5[11]) );
  FA_X1 p10_Partial_products_sum_add_23_U1_20 ( .A(p10_final_product1[26]), 
        .B(p10_final_product2_26_), .CI(
        p10_Partial_products_sum_add_23_carry_20_), .S(temp5[13]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_7 ( .A(p11_S[61]), .B(p11_C[60]), 
        .CI(p11_Partial_products_sum_add_23_carry_7_), .CO(
        p11_Partial_products_sum_add_23_carry_8_), .S(temp6[0]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_8 ( .A(p11_S[62]), .B(p11_C[61]), 
        .CI(p11_Partial_products_sum_add_23_carry_8_), .CO(
        p11_Partial_products_sum_add_23_carry_9_), .S(temp6[1]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_9 ( .A(p11_S[63]), .B(p11_C[62]), 
        .CI(p11_Partial_products_sum_add_23_carry_9_), .CO(
        p11_Partial_products_sum_add_23_carry_10_), .S(temp6[2]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_10 ( .A(p11_S[64]), .B(p11_C[63]), 
        .CI(p11_Partial_products_sum_add_23_carry_10_), .CO(
        p11_Partial_products_sum_add_23_carry_11_), .S(temp6[3]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_11 ( .A(p11_S[65]), .B(p11_C[64]), 
        .CI(p11_Partial_products_sum_add_23_carry_11_), .CO(
        p11_Partial_products_sum_add_23_carry_12_), .S(temp6[4]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_12 ( .A(p11_S[66]), .B(p11_C[65]), 
        .CI(p11_Partial_products_sum_add_23_carry_12_), .CO(
        p11_Partial_products_sum_add_23_carry_13_), .S(temp6[5]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_13 ( .A(p11_S[67]), .B(p11_C[66]), 
        .CI(p11_Partial_products_sum_add_23_carry_13_), .CO(
        p11_Partial_products_sum_add_23_carry_14_), .S(temp6[6]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_14 ( .A(p11_S[68]), .B(p11_C[67]), 
        .CI(p11_Partial_products_sum_add_23_carry_14_), .CO(
        p11_Partial_products_sum_add_23_carry_15_), .S(temp6[7]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_15 ( .A(p11_S[69]), .B(p11_C[68]), 
        .CI(p11_Partial_products_sum_add_23_carry_15_), .CO(
        p11_Partial_products_sum_add_23_carry_16_), .S(temp6[8]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_16 ( .A(p11_S[70]), .B(p11_C[69]), 
        .CI(p11_Partial_products_sum_add_23_carry_16_), .CO(
        p11_Partial_products_sum_add_23_carry_17_), .S(temp6[9]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_17 ( .A(p11_S[71]), .B(p11_C[70]), 
        .CI(p11_Partial_products_sum_add_23_carry_17_), .CO(
        p11_Partial_products_sum_add_23_carry_18_), .S(temp6[10]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_18 ( .A(p11_S[72]), .B(p11_C[71]), 
        .CI(p11_Partial_products_sum_add_23_carry_18_), .CO(
        p11_Partial_products_sum_add_23_carry_19_), .S(temp6[11]) );
  FA_X1 p11_Partial_products_sum_add_23_U1_20 ( .A(p11_final_product1[26]), 
        .B(p11_final_product2_26_), .CI(
        p11_Partial_products_sum_add_23_carry_20_), .S(temp6[13]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_7 ( .A(p9_S[61]), .B(p9_C[60]), .CI(
        p9_Partial_products_sum_add_23_carry_7_), .CO(
        p9_Partial_products_sum_add_23_carry_8_), .S(temp4[0]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_8 ( .A(p9_S[62]), .B(p9_C[61]), .CI(
        p9_Partial_products_sum_add_23_carry_8_), .CO(
        p9_Partial_products_sum_add_23_carry_9_), .S(temp4[1]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_9 ( .A(p9_S[63]), .B(p9_C[62]), .CI(
        p9_Partial_products_sum_add_23_carry_9_), .CO(
        p9_Partial_products_sum_add_23_carry_10_), .S(temp4[2]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_10 ( .A(p9_S[64]), .B(p9_C[63]), 
        .CI(p9_Partial_products_sum_add_23_carry_10_), .CO(
        p9_Partial_products_sum_add_23_carry_11_), .S(temp4[3]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_11 ( .A(p9_S[65]), .B(p9_C[64]), 
        .CI(p9_Partial_products_sum_add_23_carry_11_), .CO(
        p9_Partial_products_sum_add_23_carry_12_), .S(temp4[4]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_12 ( .A(p9_S[66]), .B(p9_C[65]), 
        .CI(p9_Partial_products_sum_add_23_carry_12_), .CO(
        p9_Partial_products_sum_add_23_carry_13_), .S(temp4[5]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_13 ( .A(p9_S[67]), .B(p9_C[66]), 
        .CI(p9_Partial_products_sum_add_23_carry_13_), .CO(
        p9_Partial_products_sum_add_23_carry_14_), .S(temp4[6]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_14 ( .A(p9_S[68]), .B(p9_C[67]), 
        .CI(p9_Partial_products_sum_add_23_carry_14_), .CO(
        p9_Partial_products_sum_add_23_carry_15_), .S(temp4[7]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_15 ( .A(p9_S[69]), .B(p9_C[68]), 
        .CI(p9_Partial_products_sum_add_23_carry_15_), .CO(
        p9_Partial_products_sum_add_23_carry_16_), .S(temp4[8]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_16 ( .A(p9_S[70]), .B(p9_C[69]), 
        .CI(p9_Partial_products_sum_add_23_carry_16_), .CO(
        p9_Partial_products_sum_add_23_carry_17_), .S(temp4[9]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_17 ( .A(p9_S[71]), .B(p9_C[70]), 
        .CI(p9_Partial_products_sum_add_23_carry_17_), .CO(
        p9_Partial_products_sum_add_23_carry_18_), .S(temp4[10]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_18 ( .A(p9_S[72]), .B(p9_C[71]), 
        .CI(p9_Partial_products_sum_add_23_carry_18_), .CO(
        p9_Partial_products_sum_add_23_carry_19_), .S(temp4[11]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_19 ( .A(p9_C[72]), .B(
        p9_final_product2_25_), .CI(p9_Partial_products_sum_add_23_carry_19_), 
        .CO(p9_Partial_products_sum_add_23_carry_20_), .S(temp4[12]) );
  FA_X1 p9_Partial_products_sum_add_23_U1_20 ( .A(p9_final_product1[26]), .B(
        p9_final_product2_26_), .CI(p9_Partial_products_sum_add_23_carry_20_), 
        .S(temp4[13]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_7 ( .A(p8_S[61]), .B(p8_C[60]), .CI(
        p8_Partial_products_sum_add_23_carry_7_), .CO(
        p8_Partial_products_sum_add_23_carry_8_), .S(temp3[0]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_8 ( .A(p8_S[62]), .B(p8_C[61]), .CI(
        p8_Partial_products_sum_add_23_carry_8_), .CO(
        p8_Partial_products_sum_add_23_carry_9_), .S(temp3[1]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_9 ( .A(p8_S[63]), .B(p8_C[62]), .CI(
        p8_Partial_products_sum_add_23_carry_9_), .CO(
        p8_Partial_products_sum_add_23_carry_10_), .S(temp3[2]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_10 ( .A(p8_S[64]), .B(p8_C[63]), 
        .CI(p8_Partial_products_sum_add_23_carry_10_), .CO(
        p8_Partial_products_sum_add_23_carry_11_), .S(temp3[3]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_11 ( .A(p8_S[65]), .B(p8_C[64]), 
        .CI(p8_Partial_products_sum_add_23_carry_11_), .CO(
        p8_Partial_products_sum_add_23_carry_12_), .S(temp3[4]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_12 ( .A(p8_S[66]), .B(p8_C[65]), 
        .CI(p8_Partial_products_sum_add_23_carry_12_), .CO(
        p8_Partial_products_sum_add_23_carry_13_), .S(temp3[5]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_13 ( .A(p8_S[67]), .B(p8_C[66]), 
        .CI(p8_Partial_products_sum_add_23_carry_13_), .CO(
        p8_Partial_products_sum_add_23_carry_14_), .S(temp3[6]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_14 ( .A(p8_S[68]), .B(p8_C[67]), 
        .CI(p8_Partial_products_sum_add_23_carry_14_), .CO(
        p8_Partial_products_sum_add_23_carry_15_), .S(temp3[7]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_15 ( .A(p8_S[69]), .B(p8_C[68]), 
        .CI(p8_Partial_products_sum_add_23_carry_15_), .CO(
        p8_Partial_products_sum_add_23_carry_16_), .S(temp3[8]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_16 ( .A(p8_S[70]), .B(p8_C[69]), 
        .CI(p8_Partial_products_sum_add_23_carry_16_), .CO(
        p8_Partial_products_sum_add_23_carry_17_), .S(temp3[9]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_17 ( .A(p8_S[71]), .B(p8_C[70]), 
        .CI(p8_Partial_products_sum_add_23_carry_17_), .CO(
        p8_Partial_products_sum_add_23_carry_18_), .S(temp3[10]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_18 ( .A(p8_S[72]), .B(p8_C[71]), 
        .CI(p8_Partial_products_sum_add_23_carry_18_), .CO(
        p8_Partial_products_sum_add_23_carry_19_), .S(temp3[11]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_19 ( .A(p8_C[72]), .B(
        p8_final_product2_25_), .CI(p8_Partial_products_sum_add_23_carry_19_), 
        .CO(p8_Partial_products_sum_add_23_carry_20_), .S(temp3[12]) );
  FA_X1 p8_Partial_products_sum_add_23_U1_20 ( .A(p8_final_product1[26]), .B(
        p8_final_product2_26_), .CI(p8_Partial_products_sum_add_23_carry_20_), 
        .S(temp3[13]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_7 ( .A(p7_S[61]), .B(p7_C[60]), .CI(
        p7_Partial_products_sum_add_23_carry_7_), .CO(
        p7_Partial_products_sum_add_23_carry_8_), .S(temp2[0]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_8 ( .A(p7_S[62]), .B(p7_C[61]), .CI(
        p7_Partial_products_sum_add_23_carry_8_), .CO(
        p7_Partial_products_sum_add_23_carry_9_), .S(temp2[1]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_9 ( .A(p7_S[63]), .B(p7_C[62]), .CI(
        p7_Partial_products_sum_add_23_carry_9_), .CO(
        p7_Partial_products_sum_add_23_carry_10_), .S(temp2[2]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_10 ( .A(p7_S[64]), .B(p7_C[63]), 
        .CI(p7_Partial_products_sum_add_23_carry_10_), .CO(
        p7_Partial_products_sum_add_23_carry_11_), .S(temp2[3]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_11 ( .A(p7_S[65]), .B(p7_C[64]), 
        .CI(p7_Partial_products_sum_add_23_carry_11_), .CO(
        p7_Partial_products_sum_add_23_carry_12_), .S(temp2[4]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_12 ( .A(p7_S[66]), .B(p7_C[65]), 
        .CI(p7_Partial_products_sum_add_23_carry_12_), .CO(
        p7_Partial_products_sum_add_23_carry_13_), .S(temp2[5]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_13 ( .A(p7_S[67]), .B(p7_C[66]), 
        .CI(p7_Partial_products_sum_add_23_carry_13_), .CO(
        p7_Partial_products_sum_add_23_carry_14_), .S(temp2[6]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_14 ( .A(p7_S[68]), .B(p7_C[67]), 
        .CI(p7_Partial_products_sum_add_23_carry_14_), .CO(
        p7_Partial_products_sum_add_23_carry_15_), .S(temp2[7]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_15 ( .A(p7_S[69]), .B(p7_C[68]), 
        .CI(p7_Partial_products_sum_add_23_carry_15_), .CO(
        p7_Partial_products_sum_add_23_carry_16_), .S(temp2[8]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_16 ( .A(p7_S[70]), .B(p7_C[69]), 
        .CI(p7_Partial_products_sum_add_23_carry_16_), .CO(
        p7_Partial_products_sum_add_23_carry_17_), .S(temp2[9]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_17 ( .A(p7_S[71]), .B(p7_C[70]), 
        .CI(p7_Partial_products_sum_add_23_carry_17_), .CO(
        p7_Partial_products_sum_add_23_carry_18_), .S(temp2[10]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_18 ( .A(p7_S[72]), .B(p7_C[71]), 
        .CI(p7_Partial_products_sum_add_23_carry_18_), .CO(
        p7_Partial_products_sum_add_23_carry_19_), .S(temp2[11]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_19 ( .A(p7_C[72]), .B(
        p7_final_product2_25_), .CI(p7_Partial_products_sum_add_23_carry_19_), 
        .CO(p7_Partial_products_sum_add_23_carry_20_), .S(temp2[12]) );
  FA_X1 p7_Partial_products_sum_add_23_U1_20 ( .A(p7_final_product1[26]), .B(
        p7_final_product2_26_), .CI(p7_Partial_products_sum_add_23_carry_20_), 
        .S(temp2[13]) );
  FA_X1 p6_Partial_products_sum_add_23_U15 ( .A(p6_S[61]), .B(p6_C[60]), .CI(
        p6_Partial_products_sum_add_23_n15), .CO(
        p6_Partial_products_sum_add_23_n14), .S(temp1[0]) );
  FA_X1 p6_Partial_products_sum_add_23_U14 ( .A(p6_S[62]), .B(p6_C[61]), .CI(
        p6_Partial_products_sum_add_23_n14), .CO(
        p6_Partial_products_sum_add_23_n13), .S(temp1[1]) );
  FA_X1 p6_Partial_products_sum_add_23_U13 ( .A(p6_S[63]), .B(p6_C[62]), .CI(
        p6_Partial_products_sum_add_23_n13), .CO(
        p6_Partial_products_sum_add_23_n12), .S(temp1[2]) );
  FA_X1 p6_Partial_products_sum_add_23_U12 ( .A(p6_S[64]), .B(p6_C[63]), .CI(
        p6_Partial_products_sum_add_23_n12), .CO(
        p6_Partial_products_sum_add_23_n11), .S(temp1[3]) );
  FA_X1 p6_Partial_products_sum_add_23_U11 ( .A(p6_S[65]), .B(p6_C[64]), .CI(
        p6_Partial_products_sum_add_23_n11), .CO(
        p6_Partial_products_sum_add_23_n10), .S(temp1[4]) );
  FA_X1 p6_Partial_products_sum_add_23_U10 ( .A(p6_S[66]), .B(p6_C[65]), .CI(
        p6_Partial_products_sum_add_23_n10), .CO(
        p6_Partial_products_sum_add_23_n9), .S(temp1[5]) );
  FA_X1 p6_Partial_products_sum_add_23_U9 ( .A(p6_S[67]), .B(p6_C[66]), .CI(
        p6_Partial_products_sum_add_23_n9), .CO(
        p6_Partial_products_sum_add_23_n8), .S(temp1[6]) );
  FA_X1 p6_Partial_products_sum_add_23_U8 ( .A(p6_S[68]), .B(p6_C[67]), .CI(
        p6_Partial_products_sum_add_23_n8), .CO(
        p6_Partial_products_sum_add_23_n7), .S(temp1[7]) );
  FA_X1 p6_Partial_products_sum_add_23_U7 ( .A(p6_S[69]), .B(p6_C[68]), .CI(
        p6_Partial_products_sum_add_23_n7), .CO(
        p6_Partial_products_sum_add_23_n6), .S(temp1[8]) );
  FA_X1 p6_Partial_products_sum_add_23_U6 ( .A(p6_S[70]), .B(p6_C[69]), .CI(
        p6_Partial_products_sum_add_23_n6), .CO(
        p6_Partial_products_sum_add_23_n5), .S(temp1[9]) );
  FA_X1 p6_Partial_products_sum_add_23_U5 ( .A(p6_S[71]), .B(p6_C[70]), .CI(
        p6_Partial_products_sum_add_23_n5), .CO(
        p6_Partial_products_sum_add_23_n4), .S(temp1[10]) );
  FA_X1 p6_Partial_products_sum_add_23_U4 ( .A(p6_S[72]), .B(p6_C[71]), .CI(
        p6_Partial_products_sum_add_23_n4), .CO(
        p6_Partial_products_sum_add_23_n3), .S(temp1[11]) );
  FA_X1 p6_Partial_products_sum_add_23_U3 ( .A(p6_C[72]), .B(
        p6_final_product2_25_), .CI(p6_Partial_products_sum_add_23_n3), .CO(
        p6_Partial_products_sum_add_23_n2), .S(temp1[12]) );
  DFFR_X2 REGISTER4_q_reg_7_ ( .D(n2502), .CK(CLK), .RN(RST_n), .Q(
        p9_Partial_products_sum_add_23_B_0_), .QN(n2801) );
  DFFR_X2 REGISTER3_q_reg_7_ ( .D(n2505), .CK(CLK), .RN(RST_n), .Q(
        p8_Partial_products_sum_add_23_B_0_), .QN(n2800) );
  DFFR_X2 REGISTER2_q_reg_7_ ( .D(n2507), .CK(CLK), .RN(RST_n), .Q(
        p7_Partial_products_sum_add_23_B_0_), .QN(n2799) );
  DFFR_X2 REGISTER1_q_reg_7_ ( .D(n2509), .CK(CLK), .RN(RST_n), .Q(
        p6_Partial_products_sum_add_23_B_0_), .QN(n2796) );
  DFFR_X1 REGISTER1_q_reg_4_ ( .D(n2533), .CK(CLK), .RN(RST_n), .Q(reg1_reg[4]), .QN(n2826) );
  DFFR_X1 REGISTER4_q_reg_6_ ( .D(n2510), .CK(CLK), .RN(RST_n), .Q(reg4_reg[6]), .QN(n2825) );
  DFFR_X1 REGISTER3_q_reg_6_ ( .D(n2513), .CK(CLK), .RN(RST_n), .Q(reg3_reg[6]), .QN(n2824) );
  DFFR_X1 REGISTER2_q_reg_6_ ( .D(n2515), .CK(CLK), .RN(RST_n), .Q(reg2_reg[6]), .QN(n2823) );
  DFFR_X1 REGISTER1_q_reg_6_ ( .D(n2517), .CK(CLK), .RN(RST_n), .Q(reg1_reg[6]), .QN(n2822) );
  AOI222_X1 U2682 ( .A1(n1384), .A2(n1385), .B1(n1384), .B2(n1382), .C1(n1385), 
        .C2(n1382), .ZN(p11_C[58]) );
  INV_X1 U2683 ( .A(B0[13]), .ZN(p6_minus_A_shifted_38_) );
  AOI21_X1 U2684 ( .B1(n2842), .B2(n1651), .A(n1640), .ZN(n1643) );
  INV_X1 U2685 ( .A(n1601), .ZN(n2621) );
  AOI22_X1 U2686 ( .A1(n1601), .A2(n1600), .B1(A1[11]), .B2(n2621), .ZN(n1378)
         );
  INV_X1 U2687 ( .A(n1941), .ZN(n2622) );
  AOI22_X1 U2688 ( .A1(n1941), .A2(n1940), .B1(A2[11]), .B2(n2622), .ZN(n1718)
         );
  INV_X1 U2689 ( .A(n83), .ZN(n2623) );
  INV_X1 U2690 ( .A(n82), .ZN(n2624) );
  AOI21_X1 U2691 ( .B1(n83), .B2(n82), .A(n80), .ZN(n2625) );
  AOI21_X1 U2692 ( .B1(n2623), .B2(n2624), .A(n2625), .ZN(n2626) );
  XNOR2_X1 U2693 ( .A(n76), .B(n78), .ZN(n2627) );
  XNOR2_X1 U2694 ( .A(n2627), .B(n79), .ZN(n2628) );
  AOI222_X1 U2695 ( .A1(p9_C[56]), .A2(n2734), .B1(p9_C[56]), .B2(p9_S[57]), 
        .C1(n2734), .C2(p9_S[57]), .ZN(n2629) );
  AOI222_X1 U2696 ( .A1(n2626), .A2(n2628), .B1(n2626), .B2(n2629), .C1(n2628), 
        .C2(n2629), .ZN(n2735) );
  INV_X1 U2697 ( .A(n409), .ZN(n2630) );
  INV_X1 U2698 ( .A(n408), .ZN(n2631) );
  AOI21_X1 U2699 ( .B1(n409), .B2(n408), .A(n406), .ZN(n2632) );
  AOI21_X1 U2700 ( .B1(n2630), .B2(n2631), .A(n2632), .ZN(n2633) );
  XNOR2_X1 U2701 ( .A(n402), .B(n404), .ZN(n2634) );
  XNOR2_X1 U2702 ( .A(n2634), .B(n405), .ZN(n2635) );
  AOI222_X1 U2703 ( .A1(p8_C[56]), .A2(n2722), .B1(p8_C[56]), .B2(p8_S[57]), 
        .C1(n2722), .C2(p8_S[57]), .ZN(n2636) );
  AOI222_X1 U2704 ( .A1(n2633), .A2(n2635), .B1(n2633), .B2(n2636), .C1(n2635), 
        .C2(n2636), .ZN(n2723) );
  AOI21_X1 U2705 ( .B1(n735), .B2(n734), .A(n732), .ZN(n2637) );
  AOI21_X1 U2706 ( .B1(n2638), .B2(n2639), .A(n2637), .ZN(n2640) );
  XNOR2_X1 U2707 ( .A(n728), .B(n730), .ZN(n2641) );
  XNOR2_X1 U2708 ( .A(n2641), .B(n731), .ZN(n2642) );
  AOI222_X1 U2709 ( .A1(p7_C[56]), .A2(n2710), .B1(p7_C[56]), .B2(p7_S[57]), 
        .C1(n2710), .C2(p7_S[57]), .ZN(n2643) );
  AOI222_X1 U2710 ( .A1(n2640), .A2(n2642), .B1(n2640), .B2(n2643), .C1(n2642), 
        .C2(n2643), .ZN(n2711) );
  INV_X1 U2711 ( .A(n735), .ZN(n2638) );
  INV_X1 U2712 ( .A(n734), .ZN(n2639) );
  XOR2_X1 U2713 ( .A(s9_add_23_DP_OP_276_9387_1_n22), .B(reg6[13]), .Z(n2644)
         );
  XNOR2_X1 U2714 ( .A(xin[13]), .B(reg7[13]), .ZN(n2645) );
  XNOR2_X1 U2715 ( .A(n2644), .B(n2645), .ZN(n2646) );
  NAND2_X1 U2716 ( .A1(s9_add_23_DP_OP_276_9387_1_n37), .A2(n2646), .ZN(n2647)
         );
  OAI211_X1 U2717 ( .C1(s9_add_23_DP_OP_276_9387_1_n37), .C2(n2646), .A(VIN), 
        .B(n2647), .ZN(n2057) );
  XOR2_X1 U2718 ( .A(A1[2]), .B(A1[1]), .Z(n3234) );
  MUX2_X1 U2719 ( .A(n3353), .B(A2[3]), .S(A2[4]), .Z(n3384) );
  MUX2_X1 U2720 ( .A(A2[6]), .B(n3385), .S(A2[5]), .Z(n3418) );
  OAI21_X1 U2721 ( .B1(n2750), .B2(p11_C[58]), .A(p11_S[59]), .ZN(n2648) );
  AND2_X1 U2722 ( .A1(n2648), .A2(n2757), .ZN(n2753) );
  OAI21_X1 U2723 ( .B1(n2770), .B2(p10_C[58]), .A(p10_S[59]), .ZN(n2649) );
  AND2_X1 U2724 ( .A1(n2649), .A2(n2777), .ZN(n2773) );
  INV_X1 U2725 ( .A(n1261), .ZN(n2650) );
  AOI22_X1 U2726 ( .A1(n1261), .A2(n1260), .B1(reg1_reg[11]), .B2(n2650), .ZN(
        n1050) );
  INV_X1 U2727 ( .A(n283), .ZN(n2651) );
  AOI22_X1 U2728 ( .A1(n283), .A2(n282), .B1(reg4_reg[11]), .B2(n2651), .ZN(
        n72) );
  INV_X1 U2729 ( .A(n609), .ZN(n2652) );
  AOI22_X1 U2730 ( .A1(n609), .A2(n608), .B1(reg3_reg[11]), .B2(n2652), .ZN(
        n398) );
  INV_X1 U2731 ( .A(n935), .ZN(n2653) );
  AOI22_X1 U2732 ( .A1(n935), .A2(n934), .B1(reg2_reg[11]), .B2(n2653), .ZN(
        n724) );
  OAI21_X1 U2733 ( .B1(p10_Partial_products_sum_add_23_carry_19_), .B2(
        p10_C[72]), .A(p10_final_product2_25_), .ZN(n2654) );
  NAND2_X1 U2734 ( .A1(n2654), .A2(n2779), .ZN(
        p10_Partial_products_sum_add_23_carry_20_) );
  OAI21_X1 U2735 ( .B1(n996), .B2(n998), .A(B0[13]), .ZN(n2655) );
  OAI21_X1 U2736 ( .B1(B0[13]), .B2(n2867), .A(n2655), .ZN(n2656) );
  XNOR2_X1 U2737 ( .A(p6_Partial_products_sum_add_23_n2), .B(n2656), .ZN(n2657) );
  XNOR2_X1 U2738 ( .A(n2657), .B(p6_final_product2_26_), .ZN(n2658) );
  INV_X1 U2739 ( .A(VIN), .ZN(n2659) );
  AOI22_X1 U2740 ( .A1(VIN), .A2(n2658), .B1(n2186), .B2(n2659), .ZN(n2447) );
  INV_X2 U2741 ( .A(A1[5]), .ZN(n3290) );
  INV_X2 U2742 ( .A(A2[5]), .ZN(n3382) );
  INV_X2 U2743 ( .A(B1[13]), .ZN(p7_minus_A_shifted_38_) );
  INV_X2 U2744 ( .A(B2[13]), .ZN(p8_minus_A_shifted_38_) );
  INV_X2 U2745 ( .A(B3[13]), .ZN(p9_minus_A_shifted_38_) );
  INV_X2 U2746 ( .A(A1[7]), .ZN(n3323) );
  INV_X2 U2747 ( .A(A2[7]), .ZN(n3415) );
  INV_X2 U2748 ( .A(B0[4]), .ZN(p6_minus_A_shifted_17_) );
  INV_X2 U2749 ( .A(B0[5]), .ZN(p6_minus_A_shifted_18_) );
  INV_X2 U2750 ( .A(B0[6]), .ZN(p6_minus_A_shifted_19_) );
  INV_X2 U2751 ( .A(B0[7]), .ZN(p6_minus_A_shifted_20_) );
  INV_X2 U2752 ( .A(B0[8]), .ZN(p6_minus_A_shifted_21_) );
  INV_X2 U2753 ( .A(B0[9]), .ZN(p6_minus_A_shifted_22_) );
  INV_X2 U2754 ( .A(B0[10]), .ZN(p6_minus_A_shifted_23_) );
  INV_X2 U2755 ( .A(B0[3]), .ZN(p6_minus_A_shifted_16_) );
  INV_X2 U2756 ( .A(B1[4]), .ZN(p7_minus_A_shifted_17_) );
  INV_X2 U2757 ( .A(B1[5]), .ZN(p7_minus_A_shifted_18_) );
  INV_X2 U2758 ( .A(B1[6]), .ZN(p7_minus_A_shifted_19_) );
  INV_X2 U2759 ( .A(B1[7]), .ZN(p7_minus_A_shifted_20_) );
  INV_X2 U2760 ( .A(B1[8]), .ZN(p7_minus_A_shifted_21_) );
  INV_X2 U2761 ( .A(B1[9]), .ZN(p7_minus_A_shifted_22_) );
  INV_X2 U2762 ( .A(B1[10]), .ZN(p7_minus_A_shifted_23_) );
  INV_X2 U2763 ( .A(B2[4]), .ZN(p8_minus_A_shifted_17_) );
  INV_X2 U2764 ( .A(B2[5]), .ZN(p8_minus_A_shifted_18_) );
  INV_X2 U2765 ( .A(B2[6]), .ZN(p8_minus_A_shifted_19_) );
  INV_X2 U2766 ( .A(B2[7]), .ZN(p8_minus_A_shifted_20_) );
  INV_X2 U2767 ( .A(B2[8]), .ZN(p8_minus_A_shifted_21_) );
  INV_X2 U2768 ( .A(B2[9]), .ZN(p8_minus_A_shifted_22_) );
  INV_X2 U2769 ( .A(B2[10]), .ZN(p8_minus_A_shifted_23_) );
  INV_X2 U2770 ( .A(B3[4]), .ZN(p9_minus_A_shifted_17_) );
  INV_X2 U2771 ( .A(B3[5]), .ZN(p9_minus_A_shifted_18_) );
  INV_X2 U2772 ( .A(B3[6]), .ZN(p9_minus_A_shifted_19_) );
  INV_X2 U2773 ( .A(B3[7]), .ZN(p9_minus_A_shifted_20_) );
  INV_X2 U2774 ( .A(B3[8]), .ZN(p9_minus_A_shifted_21_) );
  INV_X2 U2775 ( .A(B3[9]), .ZN(p9_minus_A_shifted_22_) );
  INV_X2 U2776 ( .A(B3[10]), .ZN(p9_minus_A_shifted_23_) );
  INV_X4 U2777 ( .A(VIN), .ZN(n3435) );
  INV_X1 U2778 ( .A(p10_final_product2_26_), .ZN(p10_final_product2_25_) );
  INV_X1 U2779 ( .A(p11_final_product2_26_), .ZN(p11_final_product2_25_) );
  OAI221_X1 U2780 ( .B1(reg4[11]), .B2(n1658), .C1(n2861), .C2(n1660), .A(
        n1742), .ZN(p10_C[72]) );
  OAI221_X1 U2781 ( .B1(reg2[11]), .B2(n1319), .C1(n2862), .C2(n1321), .A(
        n1402), .ZN(p11_C[72]) );
  NOR2_X2 U2782 ( .A1(A2[9]), .A2(n3433), .ZN(n1769) );
  NOR2_X2 U2783 ( .A1(A1[9]), .A2(n3432), .ZN(n1429) );
  BUF_X1 U2784 ( .A(n3234), .Z(n3260) );
  OAI21_X1 U2785 ( .B1(A2[9]), .B2(A2[10]), .A(n1744), .ZN(n1953) );
  OAI21_X1 U2786 ( .B1(A1[9]), .B2(A1[10]), .A(n1404), .ZN(n1613) );
  NAND2_X2 U2787 ( .A1(A1[8]), .A2(A1[7]), .ZN(n1421) );
  NAND2_X2 U2788 ( .A1(A2[8]), .A2(A2[7]), .ZN(n1761) );
  NOR2_X2 U2789 ( .A1(n2791), .A2(n948), .ZN(n752) );
  NOR2_X2 U2790 ( .A1(n2790), .A2(n1274), .ZN(n1078) );
  NOR2_X2 U2791 ( .A1(n2786), .A2(n622), .ZN(n426) );
  NOR2_X2 U2792 ( .A1(n1578), .A2(n1613), .ZN(n1407) );
  NOR2_X2 U2793 ( .A1(n2787), .A2(n296), .ZN(n100) );
  NOR2_X2 U2794 ( .A1(n1918), .A2(n1953), .ZN(n1747) );
  NOR2_X2 U2795 ( .A1(n2788), .A2(n654), .ZN(n447) );
  NOR2_X2 U2796 ( .A1(n2812), .A2(n980), .ZN(n773) );
  NOR2_X2 U2797 ( .A1(n2789), .A2(n328), .ZN(n121) );
  NOR2_X2 U2798 ( .A1(n2819), .A2(n1306), .ZN(n1099) );
  INV_X1 U2799 ( .A(n3120), .ZN(n2686) );
  INV_X1 U2800 ( .A(n3036), .ZN(n2687) );
  INV_X1 U2801 ( .A(n3204), .ZN(n2688) );
  INV_X1 U2802 ( .A(n2952), .ZN(n2689) );
  NOR2_X2 U2803 ( .A1(A2[11]), .A2(n1953), .ZN(n1746) );
  NOR2_X2 U2804 ( .A1(A1[11]), .A2(n1613), .ZN(n1406) );
  NOR2_X2 U2805 ( .A1(reg1_reg[11]), .A2(n1274), .ZN(n1077) );
  NOR2_X2 U2806 ( .A1(reg2_reg[11]), .A2(n948), .ZN(n751) );
  NOR2_X2 U2807 ( .A1(reg3_reg[11]), .A2(n622), .ZN(n425) );
  NOR2_X2 U2808 ( .A1(reg4_reg[11]), .A2(n296), .ZN(n99) );
  NOR2_X2 U2809 ( .A1(reg1_reg[9]), .A2(n1306), .ZN(n1098) );
  NOR2_X2 U2810 ( .A1(reg2_reg[9]), .A2(n980), .ZN(n772) );
  NOR2_X2 U2811 ( .A1(reg3_reg[9]), .A2(n654), .ZN(n446) );
  NOR2_X2 U2812 ( .A1(reg4_reg[9]), .A2(n328), .ZN(n120) );
  INV_X1 U2813 ( .A(n2924), .ZN(n2690) );
  INV_X1 U2814 ( .A(n3008), .ZN(n2691) );
  INV_X1 U2815 ( .A(n3092), .ZN(n2692) );
  INV_X1 U2816 ( .A(n3176), .ZN(n2693) );
  INV_X2 U2817 ( .A(n3415), .ZN(n3416) );
  INV_X2 U2818 ( .A(n3323), .ZN(n3324) );
  AOI222_X1 U2819 ( .A1(p6_C[54]), .A2(p6_S[55]), .B1(p6_C[54]), .B2(n2694), 
        .C1(p6_S[55]), .C2(n2694), .ZN(n2697) );
  NOR2_X1 U2820 ( .A1(p6_S[56]), .A2(p6_C[55]), .ZN(n2696) );
  NAND2_X1 U2821 ( .A1(p6_S[56]), .A2(p6_C[55]), .ZN(n2695) );
  OAI21_X1 U2822 ( .B1(n2697), .B2(n2696), .A(n2695), .ZN(n2698) );
  AOI222_X1 U2823 ( .A1(p6_C[56]), .A2(p6_S[57]), .B1(p6_C[56]), .B2(n2698), 
        .C1(p6_S[57]), .C2(n2698), .ZN(n2701) );
  NOR2_X1 U2824 ( .A1(p6_S[58]), .A2(p6_C[57]), .ZN(n2700) );
  NAND2_X1 U2825 ( .A1(p6_S[58]), .A2(p6_C[57]), .ZN(n2699) );
  OAI21_X1 U2826 ( .B1(n2701), .B2(n2700), .A(n2699), .ZN(n2702) );
  AOI222_X1 U2827 ( .A1(p6_C[58]), .A2(p6_S[59]), .B1(p6_C[58]), .B2(n2702), 
        .C1(p6_S[59]), .C2(n2702), .ZN(n2705) );
  NOR2_X1 U2828 ( .A1(p6_S[60]), .A2(p6_C[59]), .ZN(n2704) );
  NAND2_X1 U2829 ( .A1(p6_S[60]), .A2(p6_C[59]), .ZN(n2703) );
  OAI21_X1 U2830 ( .B1(n2705), .B2(n2704), .A(n2703), .ZN(
        p6_Partial_products_sum_add_23_n15) );
  AND2_X1 U2831 ( .A1(p6_S[54]), .A2(p6_Partial_products_sum_add_23_B_0_), 
        .ZN(n2694) );
  NOR2_X1 U2832 ( .A1(p7_S[56]), .A2(p7_C[55]), .ZN(n2709) );
  OAI211_X1 U2833 ( .C1(p7_S[55]), .C2(p7_C[54]), .A(
        p7_Partial_products_sum_add_23_B_0_), .B(p7_S[54]), .ZN(n2708) );
  NAND2_X1 U2834 ( .A1(p7_S[55]), .A2(p7_C[54]), .ZN(n2707) );
  NAND2_X1 U2835 ( .A1(p7_S[56]), .A2(p7_C[55]), .ZN(n2706) );
  OAI221_X1 U2836 ( .B1(n2709), .B2(n2708), .C1(n2709), .C2(n2707), .A(n2706), 
        .ZN(n2710) );
  NOR2_X1 U2837 ( .A1(p7_C[59]), .A2(p7_S[60]), .ZN(n2713) );
  NAND2_X1 U2838 ( .A1(p7_C[59]), .A2(p7_S[60]), .ZN(n2712) );
  OAI21_X1 U2839 ( .B1(n2714), .B2(n2713), .A(n2712), .ZN(
        p7_Partial_products_sum_add_23_carry_7_) );
  NAND2_X1 U2840 ( .A1(n2711), .A2(p7_C[58]), .ZN(n2715) );
  NAND2_X1 U2841 ( .A1(p7_S[59]), .A2(n2711), .ZN(n2716) );
  NAND2_X1 U2842 ( .A1(p7_S[59]), .A2(p7_C[58]), .ZN(n2717) );
  AND3_X1 U2843 ( .A1(n2717), .A2(n2716), .A3(n2715), .ZN(n2714) );
  NOR2_X1 U2844 ( .A1(p8_S[56]), .A2(p8_C[55]), .ZN(n2721) );
  OAI211_X1 U2845 ( .C1(p8_S[55]), .C2(p8_C[54]), .A(
        p8_Partial_products_sum_add_23_B_0_), .B(p8_S[54]), .ZN(n2720) );
  NAND2_X1 U2846 ( .A1(p8_S[55]), .A2(p8_C[54]), .ZN(n2719) );
  NAND2_X1 U2847 ( .A1(p8_S[56]), .A2(p8_C[55]), .ZN(n2718) );
  OAI221_X1 U2848 ( .B1(n2721), .B2(n2720), .C1(n2721), .C2(n2719), .A(n2718), 
        .ZN(n2722) );
  NOR2_X1 U2849 ( .A1(p8_C[59]), .A2(p8_S[60]), .ZN(n2725) );
  NAND2_X1 U2850 ( .A1(p8_C[59]), .A2(p8_S[60]), .ZN(n2724) );
  OAI21_X1 U2851 ( .B1(n2726), .B2(n2725), .A(n2724), .ZN(
        p8_Partial_products_sum_add_23_carry_7_) );
  NAND2_X1 U2852 ( .A1(n2723), .A2(p8_C[58]), .ZN(n2727) );
  NAND2_X1 U2853 ( .A1(p8_S[59]), .A2(n2723), .ZN(n2728) );
  NAND2_X1 U2854 ( .A1(p8_S[59]), .A2(p8_C[58]), .ZN(n2729) );
  AND3_X1 U2855 ( .A1(n2729), .A2(n2728), .A3(n2727), .ZN(n2726) );
  NOR2_X1 U2856 ( .A1(p9_S[56]), .A2(p9_C[55]), .ZN(n2733) );
  OAI211_X1 U2857 ( .C1(p9_S[55]), .C2(p9_C[54]), .A(
        p9_Partial_products_sum_add_23_B_0_), .B(p9_S[54]), .ZN(n2732) );
  NAND2_X1 U2858 ( .A1(p9_S[55]), .A2(p9_C[54]), .ZN(n2731) );
  NAND2_X1 U2859 ( .A1(p9_S[56]), .A2(p9_C[55]), .ZN(n2730) );
  OAI221_X1 U2860 ( .B1(n2733), .B2(n2732), .C1(n2733), .C2(n2731), .A(n2730), 
        .ZN(n2734) );
  NOR2_X1 U2861 ( .A1(p9_C[59]), .A2(p9_S[60]), .ZN(n2737) );
  NAND2_X1 U2862 ( .A1(p9_C[59]), .A2(p9_S[60]), .ZN(n2736) );
  OAI21_X1 U2863 ( .B1(n2738), .B2(n2737), .A(n2736), .ZN(
        p9_Partial_products_sum_add_23_carry_7_) );
  NAND2_X1 U2864 ( .A1(p9_C[58]), .A2(n2735), .ZN(n2739) );
  NAND2_X1 U2865 ( .A1(p9_S[59]), .A2(n2735), .ZN(n2740) );
  NAND2_X1 U2866 ( .A1(p9_S[59]), .A2(p9_C[58]), .ZN(n2741) );
  AND3_X1 U2867 ( .A1(n2741), .A2(n2740), .A3(n2739), .ZN(n2738) );
  NOR2_X1 U2868 ( .A1(p11_S[56]), .A2(p11_C[55]), .ZN(n2745) );
  OAI211_X1 U2869 ( .C1(p11_S[55]), .C2(p11_C[54]), .A(A1[7]), .B(p11_S[54]), 
        .ZN(n2744) );
  NAND2_X1 U2870 ( .A1(p11_S[55]), .A2(p11_C[54]), .ZN(n2743) );
  NAND2_X1 U2871 ( .A1(p11_S[56]), .A2(p11_C[55]), .ZN(n2742) );
  OAI221_X1 U2872 ( .B1(n2745), .B2(n2744), .C1(n2745), .C2(n2743), .A(n2742), 
        .ZN(n2746) );
  NOR2_X1 U2873 ( .A1(p11_S[58]), .A2(p11_C[57]), .ZN(n2748) );
  NAND2_X1 U2874 ( .A1(p11_C[57]), .A2(p11_S[58]), .ZN(n2747) );
  OAI21_X1 U2875 ( .B1(n2749), .B2(n2748), .A(n2747), .ZN(n2750) );
  NOR2_X1 U2876 ( .A1(p11_C[59]), .A2(p11_S[60]), .ZN(n2752) );
  NAND2_X1 U2877 ( .A1(p11_S[60]), .A2(p11_C[59]), .ZN(n2751) );
  OAI21_X1 U2878 ( .B1(n2753), .B2(n2752), .A(n2751), .ZN(
        p11_Partial_products_sum_add_23_carry_7_) );
  NAND2_X1 U2879 ( .A1(n2746), .A2(p11_C[56]), .ZN(n2754) );
  NAND2_X1 U2880 ( .A1(n2746), .A2(p11_S[57]), .ZN(n2755) );
  NAND2_X1 U2881 ( .A1(p11_S[57]), .A2(p11_C[56]), .ZN(n2756) );
  NAND2_X1 U2882 ( .A1(n2750), .A2(p11_C[58]), .ZN(n2757) );
  AND3_X1 U2883 ( .A1(n2756), .A2(n2755), .A3(n2754), .ZN(n2749) );
  NAND3_X1 U2884 ( .A1(n2760), .A2(n2759), .A3(n2758), .ZN(
        p11_Partial_products_sum_add_23_carry_20_) );
  NAND2_X1 U2885 ( .A1(p11_final_product2_25_), .A2(p11_C[72]), .ZN(n2758) );
  NAND2_X1 U2886 ( .A1(p11_Partial_products_sum_add_23_carry_19_), .A2(
        p11_C[72]), .ZN(n2759) );
  NAND2_X1 U2887 ( .A1(p11_Partial_products_sum_add_23_carry_19_), .A2(
        p11_final_product2_25_), .ZN(n2760) );
  XOR2_X1 U2888 ( .A(p11_Partial_products_sum_add_23_carry_19_), .B(n2761), 
        .Z(temp6[12]) );
  XOR2_X1 U2889 ( .A(p11_final_product2_25_), .B(p11_C[72]), .Z(n2761) );
  NOR2_X1 U2890 ( .A1(p10_S[56]), .A2(p10_C[55]), .ZN(n2765) );
  OAI211_X1 U2891 ( .C1(p10_S[55]), .C2(p10_C[54]), .A(A2[7]), .B(p10_S[54]), 
        .ZN(n2764) );
  NAND2_X1 U2892 ( .A1(p10_S[55]), .A2(p10_C[54]), .ZN(n2763) );
  NAND2_X1 U2893 ( .A1(p10_S[56]), .A2(p10_C[55]), .ZN(n2762) );
  OAI221_X1 U2894 ( .B1(n2765), .B2(n2764), .C1(n2778), .C2(n2763), .A(n2762), 
        .ZN(n2766) );
  NOR2_X1 U2895 ( .A1(p10_C[57]), .A2(p10_S[58]), .ZN(n2768) );
  NAND2_X1 U2896 ( .A1(p10_C[57]), .A2(p10_S[58]), .ZN(n2767) );
  OAI21_X1 U2897 ( .B1(n2769), .B2(n2768), .A(n2767), .ZN(n2770) );
  NOR2_X1 U2898 ( .A1(p10_C[59]), .A2(p10_S[60]), .ZN(n2772) );
  NAND2_X1 U2899 ( .A1(p10_C[59]), .A2(p10_S[60]), .ZN(n2771) );
  OAI21_X1 U2900 ( .B1(n2773), .B2(n2772), .A(n2771), .ZN(
        p10_Partial_products_sum_add_23_carry_7_) );
  NAND2_X1 U2901 ( .A1(n2766), .A2(p10_C[56]), .ZN(n2774) );
  NAND2_X1 U2902 ( .A1(p10_S[57]), .A2(n2766), .ZN(n2775) );
  NAND2_X1 U2903 ( .A1(p10_S[57]), .A2(p10_C[56]), .ZN(n2776) );
  NAND2_X1 U2904 ( .A1(n2770), .A2(p10_C[58]), .ZN(n2777) );
  NOR2_X1 U2905 ( .A1(p10_C[55]), .A2(p10_S[56]), .ZN(n2778) );
  AND3_X1 U2906 ( .A1(n2776), .A2(n2775), .A3(n2774), .ZN(n2769) );
  NAND2_X1 U2907 ( .A1(p10_Partial_products_sum_add_23_carry_19_), .A2(
        p10_C[72]), .ZN(n2779) );
  XOR2_X1 U2908 ( .A(p10_Partial_products_sum_add_23_carry_19_), .B(n2780), 
        .Z(temp5[12]) );
  XOR2_X1 U2909 ( .A(p10_final_product2_25_), .B(p10_C[72]), .Z(n2780) );
  NAND2_X1 U2910 ( .A1(reg7[1]), .A2(n2682), .ZN(
        s9_add_23_DP_OP_276_9387_1_n59) );
  XOR2_X1 U2911 ( .A(xin[1]), .B(reg7[1]), .Z(s9_add_23_DP_OP_276_9387_1_n60)
         );
  XOR2_X1 U2912 ( .A(mul2_reg[13]), .B(mul3_reg[13]), .Z(n2782) );
  XNOR2_X1 U2913 ( .A(mul4_reg[13]), .B(mul1_reg[13]), .ZN(n2781) );
  XNOR2_X1 U2914 ( .A(n2782), .B(n2781), .ZN(n2783) );
  XOR2_X1 U2915 ( .A(n2783), .B(s8_add_23_DP_OP_277_3998_2_n27), .Z(n2785) );
  XNOR2_X1 U2916 ( .A(s8_add_23_DP_OP_277_3998_2_n42), .B(
        s8_add_23_DP_OP_277_3998_2_n44), .ZN(n2784) );
  XNOR2_X1 U2917 ( .A(n2785), .B(n2784), .ZN(ff[13]) );
  NOR2_X2 U2918 ( .A1(n1651), .A2(n2842), .ZN(n1640) );
  INV_X2 U2919 ( .A(n3292), .ZN(n3293) );
  NOR2_X2 U2920 ( .A1(n1734), .A2(n3434), .ZN(n1770) );
  NOR2_X2 U2921 ( .A1(n1394), .A2(n1645), .ZN(n1430) );
  AOI222_X2 U2922 ( .A1(p11_muxs_out_2__7_), .A2(n1642), .B1(
        p11_muxs_out_2__7_), .B2(n1643), .C1(n1642), .C2(n1643), .ZN(n1393) );
  AOI22_X2 U2923 ( .A1(A1[4]), .A2(A1[3]), .B1(n3258), .B2(n3261), .ZN(n3262)
         );
  OR2_X1 U2924 ( .A1(VIN), .A2(n2172), .ZN(n3426) );
  AND2_X1 U2925 ( .A1(n2987), .A2(n2988), .ZN(n2855) );
  INV_X1 U2926 ( .A(B1[1]), .ZN(p7_minus_A_shifted_14_) );
  INV_X1 U2927 ( .A(B1[11]), .ZN(n2984) );
  INV_X1 U2928 ( .A(n2982), .ZN(n2983) );
  INV_X1 U2929 ( .A(n3007), .ZN(n3008) );
  INV_X1 U2930 ( .A(n3035), .ZN(n3036) );
  OR2_X1 U2931 ( .A1(VIN), .A2(n2142), .ZN(n3427) );
  AND2_X1 U2932 ( .A1(n3155), .A2(n3156), .ZN(n2857) );
  INV_X1 U2933 ( .A(B3[1]), .ZN(p9_minus_A_shifted_14_) );
  INV_X1 U2934 ( .A(B3[11]), .ZN(n3152) );
  INV_X1 U2935 ( .A(n3150), .ZN(n3151) );
  INV_X1 U2936 ( .A(n3175), .ZN(n3176) );
  INV_X1 U2937 ( .A(n3203), .ZN(n3204) );
  AND2_X1 U2938 ( .A1(n3071), .A2(n3072), .ZN(n2856) );
  INV_X1 U2939 ( .A(B2[1]), .ZN(p8_minus_A_shifted_14_) );
  INV_X1 U2940 ( .A(B2[11]), .ZN(n3068) );
  INV_X1 U2941 ( .A(n3066), .ZN(n3067) );
  INV_X1 U2942 ( .A(n3091), .ZN(n3092) );
  INV_X1 U2943 ( .A(n3119), .ZN(n3120) );
  OR2_X1 U2944 ( .A1(VIN), .A2(n2157), .ZN(n3428) );
  INV_X1 U2945 ( .A(n1065), .ZN(n1064) );
  AND2_X1 U2946 ( .A1(n2903), .A2(n2904), .ZN(n2850) );
  INV_X1 U2947 ( .A(B0[11]), .ZN(n2900) );
  INV_X1 U2948 ( .A(n2898), .ZN(n2899) );
  INV_X1 U2949 ( .A(n2923), .ZN(n2924) );
  INV_X1 U2950 ( .A(n2951), .ZN(n2952) );
  INV_X1 U2951 ( .A(n1733), .ZN(n1732) );
  AND2_X1 U2952 ( .A1(n1991), .A2(n2843), .ZN(n3422) );
  AND2_X1 U2953 ( .A1(n3333), .A2(n3334), .ZN(n2843) );
  CLKBUF_X1 U2954 ( .A(n1725), .Z(n3424) );
  INV_X1 U2955 ( .A(n1769), .ZN(n1972) );
  INV_X1 U2956 ( .A(A2[3]), .ZN(n3353) );
  INV_X1 U2957 ( .A(n1889), .ZN(n1931) );
  INV_X1 U2958 ( .A(n3330), .ZN(n3355) );
  INV_X1 U2959 ( .A(n3329), .ZN(n3330) );
  INV_X1 U2960 ( .A(A2[2]), .ZN(n3328) );
  INV_X1 U2961 ( .A(A2[1]), .ZN(n3327) );
  INV_X1 U2962 ( .A(A2[3]), .ZN(n3354) );
  INV_X1 U2963 ( .A(n3384), .ZN(n3383) );
  INV_X1 U2964 ( .A(n3418), .ZN(n3417) );
  INV_X1 U2965 ( .A(A2[6]), .ZN(n3385) );
  NAND2_X1 U2966 ( .A1(A2[9]), .A2(A2[10]), .ZN(n1744) );
  INV_X1 U2967 ( .A(n1393), .ZN(n1392) );
  AND2_X1 U2968 ( .A1(n3238), .A2(n3239), .ZN(n2842) );
  INV_X1 U2969 ( .A(n1430), .ZN(n1633) );
  INV_X1 U2970 ( .A(n1429), .ZN(n1632) );
  INV_X1 U2971 ( .A(A1[3]), .ZN(n3258) );
  INV_X1 U2972 ( .A(p11_muxs_out_2__10_), .ZN(n1614) );
  INV_X1 U2973 ( .A(n1549), .ZN(n1591) );
  INV_X1 U2974 ( .A(A1[0]), .ZN(n1657) );
  INV_X1 U2975 ( .A(n3234), .ZN(n3235) );
  INV_X1 U2976 ( .A(A1[3]), .ZN(n3259) );
  INV_X1 U2977 ( .A(n3262), .ZN(n3263) );
  INV_X1 U2978 ( .A(A1[4]), .ZN(n3261) );
  CLKBUF_X1 U2979 ( .A(n3292), .Z(n3326) );
  AOI22_X1 U2980 ( .A1(A1[6]), .A2(n3325), .B1(A1[5]), .B2(n3291), .ZN(n3292)
         );
  INV_X1 U2981 ( .A(A1[6]), .ZN(n3291) );
  INV_X1 U2982 ( .A(A1[5]), .ZN(n3325) );
  OR2_X1 U2983 ( .A1(A1[8]), .A2(A1[7]), .ZN(n3421) );
  NAND2_X1 U2984 ( .A1(A1[9]), .A2(n3431), .ZN(n1420) );
  NAND2_X1 U2985 ( .A1(A1[9]), .A2(A1[10]), .ZN(n1404) );
  AOI22_X1 U2986 ( .A1(reg2_reg[6]), .A2(n2852), .B1(reg2_reg[5]), .B2(n2823), 
        .ZN(n3035) );
  AOI22_X1 U2987 ( .A1(reg4_reg[6]), .A2(n2854), .B1(reg4_reg[5]), .B2(n2825), 
        .ZN(n3203) );
  AOI22_X1 U2988 ( .A1(reg3_reg[6]), .A2(n2853), .B1(reg3_reg[5]), .B2(n2824), 
        .ZN(n3119) );
  AOI22_X1 U2989 ( .A1(reg1_reg[6]), .A2(n2851), .B1(reg1_reg[5]), .B2(n2822), 
        .ZN(n2951) );
  NOR2_X1 U2990 ( .A1(n2866), .A2(n912), .ZN(n671) );
  NOR2_X1 U2991 ( .A1(reg2_reg[13]), .A2(n912), .ZN(n670) );
  NOR2_X1 U2992 ( .A1(n2804), .A2(n260), .ZN(n18) );
  NOR2_X1 U2993 ( .A1(reg4_reg[13]), .A2(n260), .ZN(n17) );
  NOR2_X1 U2994 ( .A1(n2805), .A2(n586), .ZN(n345) );
  NOR2_X1 U2995 ( .A1(reg3_reg[13]), .A2(n586), .ZN(n344) );
  NOR2_X1 U2996 ( .A1(n2867), .A2(n1238), .ZN(n997) );
  NOR2_X1 U2997 ( .A1(reg1_reg[13]), .A2(n1238), .ZN(n996) );
  NAND2_X1 U2998 ( .A1(n3411), .A2(n3412), .ZN(p10_muxs_out_3__19_) );
  NAND2_X1 U2999 ( .A1(n3319), .A2(n3320), .ZN(p11_muxs_out_3__19_) );
  AOI222_X1 U3000 ( .A1(p7_muxs_out_2__7_), .A2(n977), .B1(p7_muxs_out_2__7_), 
        .B2(n978), .C1(n977), .C2(n978), .ZN(n739) );
  NOR2_X1 U3001 ( .A1(n670), .A2(n672), .ZN(n3439) );
  AOI222_X1 U3002 ( .A1(p9_muxs_out_2__7_), .A2(n325), .B1(p9_muxs_out_2__7_), 
        .B2(n326), .C1(n325), .C2(n326), .ZN(n87) );
  AOI222_X1 U3003 ( .A1(n78), .A2(n79), .B1(n78), .B2(n76), .C1(n79), .C2(n76), 
        .ZN(p9_C[58]) );
  NOR2_X1 U3004 ( .A1(n17), .A2(n20), .ZN(n3437) );
  AOI222_X1 U3005 ( .A1(p8_muxs_out_2__7_), .A2(n651), .B1(p8_muxs_out_2__7_), 
        .B2(n652), .C1(n651), .C2(n652), .ZN(n413) );
  NOR2_X1 U3006 ( .A1(n344), .A2(n346), .ZN(n3438) );
  AOI222_X1 U3007 ( .A1(n1979), .A2(n1980), .B1(n1979), .B2(n1981), .C1(n1980), 
        .C2(n1981), .ZN(n1728) );
  AOI21_X1 U3008 ( .B1(n1948), .B2(n2815), .A(n1993), .ZN(n1991) );
  AOI222_X1 U3009 ( .A1(p10_muxs_out_1__8_), .A2(p10_muxs_out_2__8_), .B1(
        p10_muxs_out_1__8_), .B2(n1971), .C1(p10_muxs_out_2__8_), .C2(n1971), 
        .ZN(n1969) );
  NOR2_X1 U3010 ( .A1(n1662), .A2(n1665), .ZN(n3436) );
  AOI222_X1 U3011 ( .A1(n1639), .A2(n1640), .B1(n1641), .B2(n1639), .C1(n1640), 
        .C2(n1641), .ZN(n1388) );
  AOI21_X1 U3012 ( .B1(n1608), .B2(n2835), .A(n1653), .ZN(n1651) );
  AOI222_X1 U3013 ( .A1(n1626), .A2(n1627), .B1(n1626), .B2(n1628), .C1(n1627), 
        .C2(n1628), .ZN(n1384) );
  NAND2_X1 U3014 ( .A1(n3268), .A2(n3269), .ZN(p11_muxs_out_2__8_) );
  XOR2_X1 U3015 ( .A(n1585), .B(n1562), .Z(n1559) );
  AOI221_X1 U3016 ( .B1(n1406), .B2(reg2[9]), .C1(n1407), .C2(n2816), .A(n1458), .ZN(n1443) );
  NOR2_X1 U3017 ( .A1(n1323), .A2(n1326), .ZN(n3440) );
  AOI22_X1 U3018 ( .A1(A2[2]), .A2(A2[1]), .B1(n3327), .B2(n3328), .ZN(n3329)
         );
  AOI22_X1 U3019 ( .A1(reg1_reg[2]), .A2(reg1_reg[1]), .B1(n2864), .B2(n2792), 
        .ZN(n2898) );
  OAI221_X1 U3020 ( .B1(p6_minus_A_shifted_16_), .B2(reg1_reg[2]), .C1(B0[3]), 
        .C2(reg1_reg[3]), .A(n2899), .ZN(n2901) );
  OAI221_X1 U3021 ( .B1(reg1_reg[3]), .B2(B0[4]), .C1(n2844), .C2(
        p6_minus_A_shifted_17_), .A(n2898), .ZN(n2902) );
  NAND2_X1 U3022 ( .A1(n2901), .A2(n2902), .ZN(p6_muxs_out_1__6_) );
  OAI221_X1 U3023 ( .B1(B0[4]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_17_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2903) );
  OAI221_X1 U3024 ( .B1(reg1_reg[3]), .B2(B0[5]), .C1(n2844), .C2(
        p6_minus_A_shifted_18_), .A(n2898), .ZN(n2904) );
  OAI221_X1 U3025 ( .B1(B0[5]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_18_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2905) );
  OAI221_X1 U3026 ( .B1(reg1_reg[3]), .B2(B0[6]), .C1(n2844), .C2(
        p6_minus_A_shifted_19_), .A(n2898), .ZN(n2906) );
  NAND2_X1 U3027 ( .A1(n2905), .A2(n2906), .ZN(p6_muxs_out_1__8_) );
  OAI221_X1 U3028 ( .B1(B0[6]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_19_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2907) );
  OAI221_X1 U3029 ( .B1(reg1_reg[3]), .B2(B0[7]), .C1(n2844), .C2(
        p6_minus_A_shifted_20_), .A(n2898), .ZN(n2908) );
  NAND2_X1 U3030 ( .A1(n2907), .A2(n2908), .ZN(p6_muxs_out_1__9_) );
  OAI221_X1 U3031 ( .B1(B0[7]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_20_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2909) );
  OAI221_X1 U3032 ( .B1(reg1_reg[3]), .B2(B0[8]), .C1(n2844), .C2(
        p6_minus_A_shifted_21_), .A(n2898), .ZN(n2910) );
  NAND2_X1 U3033 ( .A1(n2909), .A2(n2910), .ZN(p6_muxs_out_1__10_) );
  OAI221_X1 U3034 ( .B1(B0[8]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_21_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2911) );
  OAI221_X1 U3035 ( .B1(reg1_reg[3]), .B2(B0[9]), .C1(n2844), .C2(
        p6_minus_A_shifted_22_), .A(n2898), .ZN(n2912) );
  NAND2_X1 U3036 ( .A1(n2911), .A2(n2912), .ZN(p6_muxs_out_1__11_) );
  OAI221_X1 U3037 ( .B1(B0[9]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_22_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2913) );
  OAI221_X1 U3038 ( .B1(reg1_reg[3]), .B2(B0[10]), .C1(n2844), .C2(
        p6_minus_A_shifted_23_), .A(n2898), .ZN(n2914) );
  NAND2_X1 U3039 ( .A1(n2913), .A2(n2914), .ZN(p6_muxs_out_1__12_) );
  OAI221_X1 U3040 ( .B1(B0[10]), .B2(reg1_reg[3]), .C1(p6_minus_A_shifted_23_), 
        .C2(reg1_reg[2]), .A(n2899), .ZN(n2915) );
  OAI221_X1 U3041 ( .B1(reg1_reg[3]), .B2(B0[11]), .C1(n2844), .C2(n2900), .A(
        n2898), .ZN(n2916) );
  NAND2_X1 U3042 ( .A1(n2915), .A2(n2916), .ZN(p6_muxs_out_1__13_) );
  OAI221_X1 U3043 ( .B1(B0[11]), .B2(reg1_reg[3]), .C1(n2900), .C2(reg1_reg[2]), .A(n2899), .ZN(n2917) );
  OAI221_X1 U3044 ( .B1(reg1_reg[3]), .B2(B0[12]), .C1(n2844), .C2(
        p6_minus_A_shifted_25_), .A(n2898), .ZN(n2918) );
  NAND2_X1 U3045 ( .A1(n2917), .A2(n2918), .ZN(p6_muxs_out_1__14_) );
  AOI22_X1 U3046 ( .A1(reg1_reg[3]), .A2(p6_minus_A_shifted_38_), .B1(B0[13]), 
        .B2(n2844), .ZN(n2919) );
  AOI22_X1 U3047 ( .A1(B0[12]), .A2(reg1_reg[2]), .B1(reg1_reg[3]), .B2(
        p6_minus_A_shifted_25_), .ZN(n2920) );
  AOI22_X1 U3048 ( .A1(n2898), .A2(n2919), .B1(n2920), .B2(n2899), .ZN(
        p6_muxs_out_1__15_) );
  AOI21_X1 U3049 ( .B1(reg1_reg[2]), .B2(reg1_reg[1]), .A(
        p6_minus_A_shifted_38_), .ZN(n2921) );
  OAI21_X1 U3050 ( .B1(reg1_reg[2]), .B2(reg1_reg[1]), .A(n2844), .ZN(n2922)
         );
  OAI22_X1 U3051 ( .A1(n2921), .A2(n2844), .B1(p6_minus_A_shifted_38_), .B2(
        n2922), .ZN(p6_muxs_out_1__16_) );
  AOI22_X1 U3052 ( .A1(reg1_reg[4]), .A2(reg1_reg[3]), .B1(n2844), .B2(n2826), 
        .ZN(n2923) );
  OAI221_X1 U3053 ( .B1(p6_minus_A_shifted_14_), .B2(reg1_reg[4]), .C1(B0[1]), 
        .C2(reg1_reg[5]), .A(n2924), .ZN(n2925) );
  OAI221_X1 U3054 ( .B1(reg1_reg[5]), .B2(B0[2]), .C1(n2851), .C2(
        p6_minus_A_shifted_15_), .A(n2923), .ZN(n2926) );
  NAND2_X1 U3055 ( .A1(n2925), .A2(n2926), .ZN(p6_muxs_out_2__6_) );
  OAI221_X1 U3056 ( .B1(B0[2]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_15_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2927) );
  OAI221_X1 U3057 ( .B1(reg1_reg[5]), .B2(B0[3]), .C1(n2851), .C2(
        p6_minus_A_shifted_16_), .A(n2923), .ZN(n2928) );
  NAND2_X1 U3058 ( .A1(n2927), .A2(n2928), .ZN(p6_muxs_out_2__7_) );
  OAI221_X1 U3059 ( .B1(B0[3]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_16_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2929) );
  OAI221_X1 U3060 ( .B1(reg1_reg[5]), .B2(B0[4]), .C1(n2851), .C2(
        p6_minus_A_shifted_17_), .A(n2923), .ZN(n2930) );
  NAND2_X1 U3061 ( .A1(n2929), .A2(n2930), .ZN(p6_muxs_out_2__8_) );
  OAI221_X1 U3062 ( .B1(B0[4]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_17_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2931) );
  OAI221_X1 U3063 ( .B1(reg1_reg[5]), .B2(B0[5]), .C1(n2851), .C2(
        p6_minus_A_shifted_18_), .A(n2923), .ZN(n2932) );
  NAND2_X1 U3064 ( .A1(n2931), .A2(n2932), .ZN(p6_muxs_out_2__9_) );
  OAI221_X1 U3065 ( .B1(B0[5]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_18_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2933) );
  OAI221_X1 U3066 ( .B1(reg1_reg[5]), .B2(B0[6]), .C1(n2851), .C2(
        p6_minus_A_shifted_19_), .A(n2923), .ZN(n2934) );
  NAND2_X1 U3067 ( .A1(n2933), .A2(n2934), .ZN(p6_muxs_out_2__10_) );
  OAI221_X1 U3068 ( .B1(B0[6]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_19_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2935) );
  OAI221_X1 U3069 ( .B1(reg1_reg[5]), .B2(B0[7]), .C1(n2851), .C2(
        p6_minus_A_shifted_20_), .A(n2923), .ZN(n2936) );
  NAND2_X1 U3070 ( .A1(n2935), .A2(n2936), .ZN(p6_muxs_out_2__11_) );
  OAI221_X1 U3071 ( .B1(B0[7]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_20_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2937) );
  OAI221_X1 U3072 ( .B1(reg1_reg[5]), .B2(B0[8]), .C1(n2851), .C2(
        p6_minus_A_shifted_21_), .A(n2923), .ZN(n2938) );
  NAND2_X1 U3073 ( .A1(n2937), .A2(n2938), .ZN(p6_muxs_out_2__12_) );
  OAI221_X1 U3074 ( .B1(B0[8]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_21_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2939) );
  OAI221_X1 U3075 ( .B1(reg1_reg[5]), .B2(B0[9]), .C1(n2851), .C2(
        p6_minus_A_shifted_22_), .A(n2923), .ZN(n2940) );
  NAND2_X1 U3076 ( .A1(n2939), .A2(n2940), .ZN(p6_muxs_out_2__13_) );
  OAI221_X1 U3077 ( .B1(B0[9]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_22_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2941) );
  OAI221_X1 U3078 ( .B1(reg1_reg[5]), .B2(B0[10]), .C1(n2851), .C2(
        p6_minus_A_shifted_23_), .A(n2923), .ZN(n2942) );
  NAND2_X1 U3079 ( .A1(n2941), .A2(n2942), .ZN(p6_muxs_out_2__14_) );
  OAI221_X1 U3080 ( .B1(B0[10]), .B2(reg1_reg[5]), .C1(p6_minus_A_shifted_23_), 
        .C2(reg1_reg[4]), .A(n2924), .ZN(n2943) );
  OAI221_X1 U3081 ( .B1(reg1_reg[5]), .B2(B0[11]), .C1(n2851), .C2(n2900), .A(
        n2923), .ZN(n2944) );
  NAND2_X1 U3082 ( .A1(n2943), .A2(n2944), .ZN(p6_muxs_out_2__15_) );
  OAI221_X1 U3083 ( .B1(B0[11]), .B2(reg1_reg[5]), .C1(n2900), .C2(reg1_reg[4]), .A(n2924), .ZN(n2945) );
  OAI221_X1 U3084 ( .B1(reg1_reg[5]), .B2(B0[12]), .C1(n2851), .C2(
        p6_minus_A_shifted_25_), .A(n2690), .ZN(n2946) );
  NAND2_X1 U3085 ( .A1(n2945), .A2(n2946), .ZN(p6_muxs_out_2__16_) );
  AOI22_X1 U3086 ( .A1(reg1_reg[5]), .A2(p6_minus_A_shifted_38_), .B1(B0[13]), 
        .B2(n2851), .ZN(n2947) );
  AOI22_X1 U3087 ( .A1(B0[12]), .A2(reg1_reg[4]), .B1(reg1_reg[5]), .B2(
        p6_minus_A_shifted_25_), .ZN(n2948) );
  AOI22_X1 U3088 ( .A1(n2690), .A2(n2947), .B1(n2948), .B2(n2924), .ZN(
        p6_muxs_out_2__17_) );
  AOI21_X1 U3089 ( .B1(reg1_reg[4]), .B2(reg1_reg[3]), .A(
        p6_minus_A_shifted_38_), .ZN(n2949) );
  OAI21_X1 U3090 ( .B1(reg1_reg[4]), .B2(reg1_reg[3]), .A(n2851), .ZN(n2950)
         );
  OAI22_X1 U3091 ( .A1(n2949), .A2(n2851), .B1(p6_minus_A_shifted_38_), .B2(
        n2950), .ZN(p6_muxs_out_2__18_) );
  NAND2_X1 U3092 ( .A1(B0[0]), .A2(n2952), .ZN(n2953) );
  XNOR2_X1 U3093 ( .A(n2953), .B(p6_Partial_products_sum_add_23_B_0_), .ZN(
        p6_muxs_out_3__6_) );
  OAI221_X1 U3094 ( .B1(B0[0]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_13_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2954) );
  OAI221_X1 U3095 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[1]), .C1(
        n2796), .C2(p6_minus_A_shifted_14_), .A(n2952), .ZN(n2955) );
  NAND2_X1 U3096 ( .A1(n2954), .A2(n2955), .ZN(p6_muxs_out_3__7_) );
  OAI221_X1 U3097 ( .B1(B0[1]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_14_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2956) );
  OAI221_X1 U3098 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[2]), .C1(
        n2796), .C2(p6_minus_A_shifted_15_), .A(n2952), .ZN(n2957) );
  NAND2_X1 U3099 ( .A1(n2956), .A2(n2957), .ZN(p6_muxs_out_3__8_) );
  OAI221_X1 U3100 ( .B1(B0[2]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_15_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2958) );
  OAI221_X1 U3101 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[3]), .C1(
        n2796), .C2(p6_minus_A_shifted_16_), .A(n2952), .ZN(n2959) );
  NAND2_X1 U3102 ( .A1(n2958), .A2(n2959), .ZN(p6_muxs_out_3__9_) );
  OAI221_X1 U3103 ( .B1(B0[3]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_16_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2960) );
  OAI221_X1 U3104 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[4]), .C1(
        n2796), .C2(p6_minus_A_shifted_17_), .A(n2952), .ZN(n2961) );
  NAND2_X1 U3105 ( .A1(n2960), .A2(n2961), .ZN(p6_muxs_out_3__10_) );
  OAI221_X1 U3106 ( .B1(B0[4]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_17_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2962) );
  OAI221_X1 U3107 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[5]), .C1(
        n2796), .C2(p6_minus_A_shifted_18_), .A(n2952), .ZN(n2963) );
  NAND2_X1 U3108 ( .A1(n2962), .A2(n2963), .ZN(p6_muxs_out_3__11_) );
  OAI221_X1 U3109 ( .B1(B0[5]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_18_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2964) );
  OAI221_X1 U3110 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[6]), .C1(
        n2796), .C2(p6_minus_A_shifted_19_), .A(n2952), .ZN(n2965) );
  NAND2_X1 U3111 ( .A1(n2964), .A2(n2965), .ZN(p6_muxs_out_3__12_) );
  OAI221_X1 U3112 ( .B1(B0[6]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_19_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2966) );
  OAI221_X1 U3113 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[7]), .C1(
        n2796), .C2(p6_minus_A_shifted_20_), .A(n2952), .ZN(n2967) );
  NAND2_X1 U3114 ( .A1(n2966), .A2(n2967), .ZN(p6_muxs_out_3__13_) );
  OAI221_X1 U3115 ( .B1(B0[7]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_20_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2968) );
  OAI221_X1 U3116 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[8]), .C1(
        n2796), .C2(p6_minus_A_shifted_21_), .A(n2952), .ZN(n2969) );
  NAND2_X1 U3117 ( .A1(n2968), .A2(n2969), .ZN(p6_muxs_out_3__14_) );
  OAI221_X1 U3118 ( .B1(B0[8]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_21_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2970) );
  OAI221_X1 U3119 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[9]), .C1(
        n2796), .C2(p6_minus_A_shifted_22_), .A(n2952), .ZN(n2971) );
  NAND2_X1 U3120 ( .A1(n2970), .A2(n2971), .ZN(p6_muxs_out_3__15_) );
  OAI221_X1 U3121 ( .B1(B0[9]), .B2(p6_Partial_products_sum_add_23_B_0_), .C1(
        p6_minus_A_shifted_22_), .C2(reg1_reg[6]), .A(n2951), .ZN(n2972) );
  OAI221_X1 U3122 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[10]), 
        .C1(n2796), .C2(p6_minus_A_shifted_23_), .A(n2952), .ZN(n2973) );
  NAND2_X1 U3123 ( .A1(n2972), .A2(n2973), .ZN(p6_muxs_out_3__16_) );
  OAI221_X1 U3124 ( .B1(B0[10]), .B2(p6_Partial_products_sum_add_23_B_0_), 
        .C1(p6_minus_A_shifted_23_), .C2(reg1_reg[6]), .A(n2689), .ZN(n2974)
         );
  OAI221_X1 U3125 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[11]), 
        .C1(n2796), .C2(n2900), .A(n2952), .ZN(n2975) );
  NAND2_X1 U3126 ( .A1(n2974), .A2(n2975), .ZN(p6_muxs_out_3__17_) );
  OAI221_X1 U3127 ( .B1(B0[11]), .B2(p6_Partial_products_sum_add_23_B_0_), 
        .C1(n2900), .C2(reg1_reg[6]), .A(n2689), .ZN(n2976) );
  OAI221_X1 U3128 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[12]), 
        .C1(n2796), .C2(p6_minus_A_shifted_25_), .A(n2952), .ZN(n2977) );
  NAND2_X1 U3129 ( .A1(n2976), .A2(n2977), .ZN(p6_muxs_out_3__18_) );
  OAI221_X1 U3130 ( .B1(B0[12]), .B2(p6_Partial_products_sum_add_23_B_0_), 
        .C1(p6_minus_A_shifted_25_), .C2(reg1_reg[6]), .A(n2689), .ZN(n2978)
         );
  OAI221_X1 U3131 ( .B1(p6_Partial_products_sum_add_23_B_0_), .B2(B0[13]), 
        .C1(n2796), .C2(p6_minus_A_shifted_38_), .A(n2952), .ZN(n2979) );
  NAND2_X1 U3132 ( .A1(n2978), .A2(n2979), .ZN(p6_muxs_out_3__19_) );
  AOI21_X1 U3133 ( .B1(reg1_reg[6]), .B2(reg1_reg[5]), .A(
        p6_minus_A_shifted_38_), .ZN(n2980) );
  OAI21_X1 U3134 ( .B1(reg1_reg[6]), .B2(reg1_reg[5]), .A(n2796), .ZN(n2981)
         );
  OAI22_X1 U3135 ( .A1(n2980), .A2(n2796), .B1(p6_minus_A_shifted_38_), .B2(
        n2981), .ZN(p6_muxs_out_3__20_) );
  AOI22_X1 U3136 ( .A1(reg2_reg[2]), .A2(reg2_reg[1]), .B1(n2865), .B2(n2793), 
        .ZN(n2982) );
  OAI221_X1 U3137 ( .B1(p7_minus_A_shifted_16_), .B2(reg2_reg[2]), .C1(B1[3]), 
        .C2(reg2_reg[3]), .A(n2983), .ZN(n2985) );
  OAI221_X1 U3138 ( .B1(reg2_reg[3]), .B2(B1[4]), .C1(n2845), .C2(
        p7_minus_A_shifted_17_), .A(n2982), .ZN(n2986) );
  NAND2_X1 U3139 ( .A1(n2985), .A2(n2986), .ZN(p7_muxs_out_1__6_) );
  OAI221_X1 U3140 ( .B1(B1[4]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_17_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2987) );
  OAI221_X1 U3141 ( .B1(reg2_reg[3]), .B2(B1[5]), .C1(n2845), .C2(
        p7_minus_A_shifted_18_), .A(n2982), .ZN(n2988) );
  OAI221_X1 U3142 ( .B1(B1[5]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_18_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2989) );
  OAI221_X1 U3143 ( .B1(reg2_reg[3]), .B2(B1[6]), .C1(n2845), .C2(
        p7_minus_A_shifted_19_), .A(n2982), .ZN(n2990) );
  NAND2_X1 U3144 ( .A1(n2989), .A2(n2990), .ZN(p7_muxs_out_1__8_) );
  OAI221_X1 U3145 ( .B1(B1[6]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_19_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2991) );
  OAI221_X1 U3146 ( .B1(reg2_reg[3]), .B2(B1[7]), .C1(n2845), .C2(
        p7_minus_A_shifted_20_), .A(n2982), .ZN(n2992) );
  NAND2_X1 U3147 ( .A1(n2991), .A2(n2992), .ZN(p7_muxs_out_1__9_) );
  OAI221_X1 U3148 ( .B1(B1[7]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_20_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2993) );
  OAI221_X1 U3149 ( .B1(reg2_reg[3]), .B2(B1[8]), .C1(n2845), .C2(
        p7_minus_A_shifted_21_), .A(n2982), .ZN(n2994) );
  NAND2_X1 U3150 ( .A1(n2993), .A2(n2994), .ZN(p7_muxs_out_1__10_) );
  OAI221_X1 U3151 ( .B1(B1[8]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_21_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2995) );
  OAI221_X1 U3152 ( .B1(reg2_reg[3]), .B2(B1[9]), .C1(n2845), .C2(
        p7_minus_A_shifted_22_), .A(n2982), .ZN(n2996) );
  NAND2_X1 U3153 ( .A1(n2995), .A2(n2996), .ZN(p7_muxs_out_1__11_) );
  OAI221_X1 U3154 ( .B1(B1[9]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_22_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2997) );
  OAI221_X1 U3155 ( .B1(reg2_reg[3]), .B2(B1[10]), .C1(n2845), .C2(
        p7_minus_A_shifted_23_), .A(n2982), .ZN(n2998) );
  NAND2_X1 U3156 ( .A1(n2997), .A2(n2998), .ZN(p7_muxs_out_1__12_) );
  OAI221_X1 U3157 ( .B1(B1[10]), .B2(reg2_reg[3]), .C1(p7_minus_A_shifted_23_), 
        .C2(reg2_reg[2]), .A(n2983), .ZN(n2999) );
  OAI221_X1 U3158 ( .B1(reg2_reg[3]), .B2(B1[11]), .C1(n2845), .C2(n2984), .A(
        n2982), .ZN(n3000) );
  NAND2_X1 U3159 ( .A1(n2999), .A2(n3000), .ZN(p7_muxs_out_1__13_) );
  OAI221_X1 U3160 ( .B1(B1[11]), .B2(reg2_reg[3]), .C1(n2984), .C2(reg2_reg[2]), .A(n2983), .ZN(n3001) );
  OAI221_X1 U3161 ( .B1(reg2_reg[3]), .B2(B1[12]), .C1(n2845), .C2(
        p7_minus_A_shifted_25_), .A(n2982), .ZN(n3002) );
  NAND2_X1 U3162 ( .A1(n3001), .A2(n3002), .ZN(p7_muxs_out_1__14_) );
  AOI22_X1 U3163 ( .A1(reg2_reg[3]), .A2(p7_minus_A_shifted_38_), .B1(B1[13]), 
        .B2(n2845), .ZN(n3003) );
  AOI22_X1 U3164 ( .A1(B1[12]), .A2(reg2_reg[2]), .B1(reg2_reg[3]), .B2(
        p7_minus_A_shifted_25_), .ZN(n3004) );
  AOI22_X1 U3165 ( .A1(n2982), .A2(n3003), .B1(n3004), .B2(n2983), .ZN(
        p7_muxs_out_1__15_) );
  AOI21_X1 U3166 ( .B1(reg2_reg[2]), .B2(reg2_reg[1]), .A(
        p7_minus_A_shifted_38_), .ZN(n3005) );
  OAI21_X1 U3167 ( .B1(reg2_reg[2]), .B2(reg2_reg[1]), .A(n2845), .ZN(n3006)
         );
  OAI22_X1 U3168 ( .A1(n3005), .A2(n2845), .B1(p7_minus_A_shifted_38_), .B2(
        n3006), .ZN(p7_muxs_out_1__16_) );
  AOI22_X1 U3169 ( .A1(reg2_reg[4]), .A2(reg2_reg[3]), .B1(n2845), .B2(n2827), 
        .ZN(n3007) );
  OAI221_X1 U3170 ( .B1(p7_minus_A_shifted_14_), .B2(reg2_reg[4]), .C1(B1[1]), 
        .C2(reg2_reg[5]), .A(n3008), .ZN(n3009) );
  OAI221_X1 U3171 ( .B1(reg2_reg[5]), .B2(B1[2]), .C1(n2852), .C2(
        p7_minus_A_shifted_15_), .A(n3007), .ZN(n3010) );
  NAND2_X1 U3172 ( .A1(n3009), .A2(n3010), .ZN(p7_muxs_out_2__6_) );
  OAI221_X1 U3173 ( .B1(B1[2]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_15_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3011) );
  OAI221_X1 U3174 ( .B1(reg2_reg[5]), .B2(B1[3]), .C1(n2852), .C2(
        p7_minus_A_shifted_16_), .A(n3007), .ZN(n3012) );
  NAND2_X1 U3175 ( .A1(n3011), .A2(n3012), .ZN(p7_muxs_out_2__7_) );
  OAI221_X1 U3176 ( .B1(B1[3]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_16_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3013) );
  OAI221_X1 U3177 ( .B1(reg2_reg[5]), .B2(B1[4]), .C1(n2852), .C2(
        p7_minus_A_shifted_17_), .A(n3007), .ZN(n3014) );
  NAND2_X1 U3178 ( .A1(n3013), .A2(n3014), .ZN(p7_muxs_out_2__8_) );
  OAI221_X1 U3179 ( .B1(B1[4]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_17_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3015) );
  OAI221_X1 U3180 ( .B1(reg2_reg[5]), .B2(B1[5]), .C1(n2852), .C2(
        p7_minus_A_shifted_18_), .A(n3007), .ZN(n3016) );
  NAND2_X1 U3181 ( .A1(n3015), .A2(n3016), .ZN(p7_muxs_out_2__9_) );
  OAI221_X1 U3182 ( .B1(B1[5]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_18_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3017) );
  OAI221_X1 U3183 ( .B1(reg2_reg[5]), .B2(B1[6]), .C1(n2852), .C2(
        p7_minus_A_shifted_19_), .A(n3007), .ZN(n3018) );
  NAND2_X1 U3184 ( .A1(n3017), .A2(n3018), .ZN(p7_muxs_out_2__10_) );
  OAI221_X1 U3185 ( .B1(B1[6]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_19_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3019) );
  OAI221_X1 U3186 ( .B1(reg2_reg[5]), .B2(B1[7]), .C1(n2852), .C2(
        p7_minus_A_shifted_20_), .A(n3007), .ZN(n3020) );
  NAND2_X1 U3187 ( .A1(n3019), .A2(n3020), .ZN(p7_muxs_out_2__11_) );
  OAI221_X1 U3188 ( .B1(B1[7]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_20_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3021) );
  OAI221_X1 U3189 ( .B1(reg2_reg[5]), .B2(B1[8]), .C1(n2852), .C2(
        p7_minus_A_shifted_21_), .A(n3007), .ZN(n3022) );
  NAND2_X1 U3190 ( .A1(n3021), .A2(n3022), .ZN(p7_muxs_out_2__12_) );
  OAI221_X1 U3191 ( .B1(B1[8]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_21_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3023) );
  OAI221_X1 U3192 ( .B1(reg2_reg[5]), .B2(B1[9]), .C1(n2852), .C2(
        p7_minus_A_shifted_22_), .A(n3007), .ZN(n3024) );
  NAND2_X1 U3193 ( .A1(n3023), .A2(n3024), .ZN(p7_muxs_out_2__13_) );
  OAI221_X1 U3194 ( .B1(B1[9]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_22_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3025) );
  OAI221_X1 U3195 ( .B1(reg2_reg[5]), .B2(B1[10]), .C1(n2852), .C2(
        p7_minus_A_shifted_23_), .A(n3007), .ZN(n3026) );
  NAND2_X1 U3196 ( .A1(n3025), .A2(n3026), .ZN(p7_muxs_out_2__14_) );
  OAI221_X1 U3197 ( .B1(B1[10]), .B2(reg2_reg[5]), .C1(p7_minus_A_shifted_23_), 
        .C2(reg2_reg[4]), .A(n3008), .ZN(n3027) );
  OAI221_X1 U3198 ( .B1(reg2_reg[5]), .B2(B1[11]), .C1(n2852), .C2(n2984), .A(
        n3007), .ZN(n3028) );
  NAND2_X1 U3199 ( .A1(n3027), .A2(n3028), .ZN(p7_muxs_out_2__15_) );
  OAI221_X1 U3200 ( .B1(B1[11]), .B2(reg2_reg[5]), .C1(n2984), .C2(reg2_reg[4]), .A(n3008), .ZN(n3029) );
  OAI221_X1 U3201 ( .B1(reg2_reg[5]), .B2(B1[12]), .C1(n2852), .C2(
        p7_minus_A_shifted_25_), .A(n2691), .ZN(n3030) );
  NAND2_X1 U3202 ( .A1(n3029), .A2(n3030), .ZN(p7_muxs_out_2__16_) );
  AOI22_X1 U3203 ( .A1(reg2_reg[5]), .A2(p7_minus_A_shifted_38_), .B1(B1[13]), 
        .B2(n2852), .ZN(n3031) );
  AOI22_X1 U3204 ( .A1(B1[12]), .A2(reg2_reg[4]), .B1(reg2_reg[5]), .B2(
        p7_minus_A_shifted_25_), .ZN(n3032) );
  AOI22_X1 U3205 ( .A1(n2691), .A2(n3031), .B1(n3032), .B2(n3008), .ZN(
        p7_muxs_out_2__17_) );
  AOI21_X1 U3206 ( .B1(reg2_reg[4]), .B2(reg2_reg[3]), .A(
        p7_minus_A_shifted_38_), .ZN(n3033) );
  OAI21_X1 U3207 ( .B1(reg2_reg[4]), .B2(reg2_reg[3]), .A(n2852), .ZN(n3034)
         );
  OAI22_X1 U3208 ( .A1(n3033), .A2(n2852), .B1(p7_minus_A_shifted_38_), .B2(
        n3034), .ZN(p7_muxs_out_2__18_) );
  NAND2_X1 U3209 ( .A1(B1[0]), .A2(n3036), .ZN(n3037) );
  XNOR2_X1 U3210 ( .A(n3037), .B(p7_Partial_products_sum_add_23_B_0_), .ZN(
        p7_muxs_out_3__6_) );
  OAI221_X1 U3211 ( .B1(B1[0]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_13_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3038) );
  OAI221_X1 U3212 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[1]), .C1(
        n2799), .C2(p7_minus_A_shifted_14_), .A(n3036), .ZN(n3039) );
  NAND2_X1 U3213 ( .A1(n3038), .A2(n3039), .ZN(p7_muxs_out_3__7_) );
  OAI221_X1 U3214 ( .B1(B1[1]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_14_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3040) );
  OAI221_X1 U3215 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[2]), .C1(
        n2799), .C2(p7_minus_A_shifted_15_), .A(n3036), .ZN(n3041) );
  NAND2_X1 U3216 ( .A1(n3040), .A2(n3041), .ZN(p7_muxs_out_3__8_) );
  OAI221_X1 U3217 ( .B1(B1[2]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_15_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3042) );
  OAI221_X1 U3218 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[3]), .C1(
        n2799), .C2(p7_minus_A_shifted_16_), .A(n3036), .ZN(n3043) );
  NAND2_X1 U3219 ( .A1(n3042), .A2(n3043), .ZN(p7_muxs_out_3__9_) );
  OAI221_X1 U3220 ( .B1(B1[3]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_16_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3044) );
  OAI221_X1 U3221 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[4]), .C1(
        n2799), .C2(p7_minus_A_shifted_17_), .A(n3036), .ZN(n3045) );
  NAND2_X1 U3222 ( .A1(n3044), .A2(n3045), .ZN(p7_muxs_out_3__10_) );
  OAI221_X1 U3223 ( .B1(B1[4]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_17_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3046) );
  OAI221_X1 U3224 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[5]), .C1(
        n2799), .C2(p7_minus_A_shifted_18_), .A(n3036), .ZN(n3047) );
  NAND2_X1 U3225 ( .A1(n3046), .A2(n3047), .ZN(p7_muxs_out_3__11_) );
  OAI221_X1 U3226 ( .B1(B1[5]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_18_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3048) );
  OAI221_X1 U3227 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[6]), .C1(
        n2799), .C2(p7_minus_A_shifted_19_), .A(n3036), .ZN(n3049) );
  NAND2_X1 U3228 ( .A1(n3048), .A2(n3049), .ZN(p7_muxs_out_3__12_) );
  OAI221_X1 U3229 ( .B1(B1[6]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_19_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3050) );
  OAI221_X1 U3230 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[7]), .C1(
        n2799), .C2(p7_minus_A_shifted_20_), .A(n3036), .ZN(n3051) );
  NAND2_X1 U3231 ( .A1(n3050), .A2(n3051), .ZN(p7_muxs_out_3__13_) );
  OAI221_X1 U3232 ( .B1(B1[7]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_20_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3052) );
  OAI221_X1 U3233 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[8]), .C1(
        n2799), .C2(p7_minus_A_shifted_21_), .A(n3036), .ZN(n3053) );
  NAND2_X1 U3234 ( .A1(n3052), .A2(n3053), .ZN(p7_muxs_out_3__14_) );
  OAI221_X1 U3235 ( .B1(B1[8]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_21_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3054) );
  OAI221_X1 U3236 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[9]), .C1(
        n2799), .C2(p7_minus_A_shifted_22_), .A(n3036), .ZN(n3055) );
  NAND2_X1 U3237 ( .A1(n3054), .A2(n3055), .ZN(p7_muxs_out_3__15_) );
  OAI221_X1 U3238 ( .B1(B1[9]), .B2(p7_Partial_products_sum_add_23_B_0_), .C1(
        p7_minus_A_shifted_22_), .C2(reg2_reg[6]), .A(n3035), .ZN(n3056) );
  OAI221_X1 U3239 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[10]), 
        .C1(n2799), .C2(p7_minus_A_shifted_23_), .A(n3036), .ZN(n3057) );
  NAND2_X1 U3240 ( .A1(n3056), .A2(n3057), .ZN(p7_muxs_out_3__16_) );
  OAI221_X1 U3241 ( .B1(B1[10]), .B2(p7_Partial_products_sum_add_23_B_0_), 
        .C1(p7_minus_A_shifted_23_), .C2(reg2_reg[6]), .A(n2687), .ZN(n3058)
         );
  OAI221_X1 U3242 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[11]), 
        .C1(n2799), .C2(n2984), .A(n3036), .ZN(n3059) );
  NAND2_X1 U3243 ( .A1(n3058), .A2(n3059), .ZN(p7_muxs_out_3__17_) );
  OAI221_X1 U3244 ( .B1(B1[11]), .B2(p7_Partial_products_sum_add_23_B_0_), 
        .C1(n2984), .C2(reg2_reg[6]), .A(n2687), .ZN(n3060) );
  OAI221_X1 U3245 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[12]), 
        .C1(n2799), .C2(p7_minus_A_shifted_25_), .A(n3036), .ZN(n3061) );
  NAND2_X1 U3246 ( .A1(n3060), .A2(n3061), .ZN(p7_muxs_out_3__18_) );
  OAI221_X1 U3247 ( .B1(B1[12]), .B2(p7_Partial_products_sum_add_23_B_0_), 
        .C1(p7_minus_A_shifted_25_), .C2(reg2_reg[6]), .A(n2687), .ZN(n3062)
         );
  OAI221_X1 U3248 ( .B1(p7_Partial_products_sum_add_23_B_0_), .B2(B1[13]), 
        .C1(n2799), .C2(p7_minus_A_shifted_38_), .A(n3036), .ZN(n3063) );
  NAND2_X1 U3249 ( .A1(n3062), .A2(n3063), .ZN(p7_muxs_out_3__19_) );
  AOI21_X1 U3250 ( .B1(reg2_reg[6]), .B2(reg2_reg[5]), .A(
        p7_minus_A_shifted_38_), .ZN(n3064) );
  OAI21_X1 U3251 ( .B1(reg2_reg[6]), .B2(reg2_reg[5]), .A(n2799), .ZN(n3065)
         );
  OAI22_X1 U3252 ( .A1(n3064), .A2(n2799), .B1(p7_minus_A_shifted_38_), .B2(
        n3065), .ZN(p7_muxs_out_3__20_) );
  AOI22_X1 U3253 ( .A1(reg3_reg[2]), .A2(reg3_reg[1]), .B1(n2840), .B2(n2794), 
        .ZN(n3066) );
  OAI221_X1 U3254 ( .B1(p8_minus_A_shifted_16_), .B2(reg3_reg[2]), .C1(B2[3]), 
        .C2(reg3_reg[3]), .A(n3067), .ZN(n3069) );
  OAI221_X1 U3255 ( .B1(reg3_reg[3]), .B2(B2[4]), .C1(n2846), .C2(
        p8_minus_A_shifted_17_), .A(n3066), .ZN(n3070) );
  NAND2_X1 U3256 ( .A1(n3069), .A2(n3070), .ZN(p8_muxs_out_1__6_) );
  OAI221_X1 U3257 ( .B1(B2[4]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_17_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3071) );
  OAI221_X1 U3258 ( .B1(reg3_reg[3]), .B2(B2[5]), .C1(n2846), .C2(
        p8_minus_A_shifted_18_), .A(n3066), .ZN(n3072) );
  OAI221_X1 U3259 ( .B1(B2[5]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_18_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3073) );
  OAI221_X1 U3260 ( .B1(reg3_reg[3]), .B2(B2[6]), .C1(n2846), .C2(
        p8_minus_A_shifted_19_), .A(n3066), .ZN(n3074) );
  NAND2_X1 U3261 ( .A1(n3073), .A2(n3074), .ZN(p8_muxs_out_1__8_) );
  OAI221_X1 U3262 ( .B1(B2[6]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_19_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3075) );
  OAI221_X1 U3263 ( .B1(reg3_reg[3]), .B2(B2[7]), .C1(n2846), .C2(
        p8_minus_A_shifted_20_), .A(n3066), .ZN(n3076) );
  NAND2_X1 U3264 ( .A1(n3075), .A2(n3076), .ZN(p8_muxs_out_1__9_) );
  OAI221_X1 U3265 ( .B1(B2[7]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_20_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3077) );
  OAI221_X1 U3266 ( .B1(reg3_reg[3]), .B2(B2[8]), .C1(n2846), .C2(
        p8_minus_A_shifted_21_), .A(n3066), .ZN(n3078) );
  NAND2_X1 U3267 ( .A1(n3077), .A2(n3078), .ZN(p8_muxs_out_1__10_) );
  OAI221_X1 U3268 ( .B1(B2[8]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_21_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3079) );
  OAI221_X1 U3269 ( .B1(reg3_reg[3]), .B2(B2[9]), .C1(n2846), .C2(
        p8_minus_A_shifted_22_), .A(n3066), .ZN(n3080) );
  NAND2_X1 U3270 ( .A1(n3079), .A2(n3080), .ZN(p8_muxs_out_1__11_) );
  OAI221_X1 U3271 ( .B1(B2[9]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_22_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3081) );
  OAI221_X1 U3272 ( .B1(reg3_reg[3]), .B2(B2[10]), .C1(n2846), .C2(
        p8_minus_A_shifted_23_), .A(n3066), .ZN(n3082) );
  NAND2_X1 U3273 ( .A1(n3081), .A2(n3082), .ZN(p8_muxs_out_1__12_) );
  OAI221_X1 U3274 ( .B1(B2[10]), .B2(reg3_reg[3]), .C1(p8_minus_A_shifted_23_), 
        .C2(reg3_reg[2]), .A(n3067), .ZN(n3083) );
  OAI221_X1 U3275 ( .B1(reg3_reg[3]), .B2(B2[11]), .C1(n2846), .C2(n3068), .A(
        n3066), .ZN(n3084) );
  NAND2_X1 U3276 ( .A1(n3083), .A2(n3084), .ZN(p8_muxs_out_1__13_) );
  OAI221_X1 U3277 ( .B1(B2[11]), .B2(reg3_reg[3]), .C1(n3068), .C2(reg3_reg[2]), .A(n3067), .ZN(n3085) );
  OAI221_X1 U3278 ( .B1(reg3_reg[3]), .B2(B2[12]), .C1(n2846), .C2(
        p8_minus_A_shifted_25_), .A(n3066), .ZN(n3086) );
  NAND2_X1 U3279 ( .A1(n3085), .A2(n3086), .ZN(p8_muxs_out_1__14_) );
  AOI22_X1 U3280 ( .A1(reg3_reg[3]), .A2(p8_minus_A_shifted_38_), .B1(B2[13]), 
        .B2(n2846), .ZN(n3087) );
  AOI22_X1 U3281 ( .A1(B2[12]), .A2(reg3_reg[2]), .B1(reg3_reg[3]), .B2(
        p8_minus_A_shifted_25_), .ZN(n3088) );
  AOI22_X1 U3282 ( .A1(n3066), .A2(n3087), .B1(n3088), .B2(n3067), .ZN(
        p8_muxs_out_1__15_) );
  AOI21_X1 U3283 ( .B1(reg3_reg[2]), .B2(reg3_reg[1]), .A(
        p8_minus_A_shifted_38_), .ZN(n3089) );
  OAI21_X1 U3284 ( .B1(reg3_reg[2]), .B2(reg3_reg[1]), .A(n2846), .ZN(n3090)
         );
  OAI22_X1 U3285 ( .A1(n3089), .A2(n2846), .B1(p8_minus_A_shifted_38_), .B2(
        n3090), .ZN(p8_muxs_out_1__16_) );
  AOI22_X1 U3286 ( .A1(reg3_reg[4]), .A2(reg3_reg[3]), .B1(n2846), .B2(n2828), 
        .ZN(n3091) );
  OAI221_X1 U3287 ( .B1(p8_minus_A_shifted_14_), .B2(reg3_reg[4]), .C1(B2[1]), 
        .C2(reg3_reg[5]), .A(n3092), .ZN(n3093) );
  OAI221_X1 U3288 ( .B1(reg3_reg[5]), .B2(B2[2]), .C1(n2853), .C2(
        p8_minus_A_shifted_15_), .A(n3091), .ZN(n3094) );
  NAND2_X1 U3289 ( .A1(n3093), .A2(n3094), .ZN(p8_muxs_out_2__6_) );
  OAI221_X1 U3290 ( .B1(B2[2]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_15_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3095) );
  OAI221_X1 U3291 ( .B1(reg3_reg[5]), .B2(B2[3]), .C1(n2853), .C2(
        p8_minus_A_shifted_16_), .A(n3091), .ZN(n3096) );
  NAND2_X1 U3292 ( .A1(n3095), .A2(n3096), .ZN(p8_muxs_out_2__7_) );
  OAI221_X1 U3293 ( .B1(B2[3]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_16_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3097) );
  OAI221_X1 U3294 ( .B1(reg3_reg[5]), .B2(B2[4]), .C1(n2853), .C2(
        p8_minus_A_shifted_17_), .A(n3091), .ZN(n3098) );
  NAND2_X1 U3295 ( .A1(n3097), .A2(n3098), .ZN(p8_muxs_out_2__8_) );
  OAI221_X1 U3296 ( .B1(B2[4]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_17_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3099) );
  OAI221_X1 U3297 ( .B1(reg3_reg[5]), .B2(B2[5]), .C1(n2853), .C2(
        p8_minus_A_shifted_18_), .A(n3091), .ZN(n3100) );
  NAND2_X1 U3298 ( .A1(n3099), .A2(n3100), .ZN(p8_muxs_out_2__9_) );
  OAI221_X1 U3299 ( .B1(B2[5]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_18_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3101) );
  OAI221_X1 U3300 ( .B1(reg3_reg[5]), .B2(B2[6]), .C1(n2853), .C2(
        p8_minus_A_shifted_19_), .A(n3091), .ZN(n3102) );
  NAND2_X1 U3301 ( .A1(n3101), .A2(n3102), .ZN(p8_muxs_out_2__10_) );
  OAI221_X1 U3302 ( .B1(B2[6]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_19_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3103) );
  OAI221_X1 U3303 ( .B1(reg3_reg[5]), .B2(B2[7]), .C1(n2853), .C2(
        p8_minus_A_shifted_20_), .A(n3091), .ZN(n3104) );
  NAND2_X1 U3304 ( .A1(n3103), .A2(n3104), .ZN(p8_muxs_out_2__11_) );
  OAI221_X1 U3305 ( .B1(B2[7]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_20_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3105) );
  OAI221_X1 U3306 ( .B1(reg3_reg[5]), .B2(B2[8]), .C1(n2853), .C2(
        p8_minus_A_shifted_21_), .A(n3091), .ZN(n3106) );
  NAND2_X1 U3307 ( .A1(n3105), .A2(n3106), .ZN(p8_muxs_out_2__12_) );
  OAI221_X1 U3308 ( .B1(B2[8]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_21_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3107) );
  OAI221_X1 U3309 ( .B1(reg3_reg[5]), .B2(B2[9]), .C1(n2853), .C2(
        p8_minus_A_shifted_22_), .A(n3091), .ZN(n3108) );
  NAND2_X1 U3310 ( .A1(n3107), .A2(n3108), .ZN(p8_muxs_out_2__13_) );
  OAI221_X1 U3311 ( .B1(B2[9]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_22_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3109) );
  OAI221_X1 U3312 ( .B1(reg3_reg[5]), .B2(B2[10]), .C1(n2853), .C2(
        p8_minus_A_shifted_23_), .A(n3091), .ZN(n3110) );
  NAND2_X1 U3313 ( .A1(n3109), .A2(n3110), .ZN(p8_muxs_out_2__14_) );
  OAI221_X1 U3314 ( .B1(B2[10]), .B2(reg3_reg[5]), .C1(p8_minus_A_shifted_23_), 
        .C2(reg3_reg[4]), .A(n3092), .ZN(n3111) );
  OAI221_X1 U3315 ( .B1(reg3_reg[5]), .B2(B2[11]), .C1(n2853), .C2(n3068), .A(
        n3091), .ZN(n3112) );
  NAND2_X1 U3316 ( .A1(n3111), .A2(n3112), .ZN(p8_muxs_out_2__15_) );
  OAI221_X1 U3317 ( .B1(B2[11]), .B2(reg3_reg[5]), .C1(n3068), .C2(reg3_reg[4]), .A(n3092), .ZN(n3113) );
  OAI221_X1 U3318 ( .B1(reg3_reg[5]), .B2(B2[12]), .C1(n2853), .C2(
        p8_minus_A_shifted_25_), .A(n2692), .ZN(n3114) );
  NAND2_X1 U3319 ( .A1(n3113), .A2(n3114), .ZN(p8_muxs_out_2__16_) );
  AOI22_X1 U3320 ( .A1(reg3_reg[5]), .A2(p8_minus_A_shifted_38_), .B1(B2[13]), 
        .B2(n2853), .ZN(n3115) );
  AOI22_X1 U3321 ( .A1(B2[12]), .A2(reg3_reg[4]), .B1(reg3_reg[5]), .B2(
        p8_minus_A_shifted_25_), .ZN(n3116) );
  AOI22_X1 U3322 ( .A1(n2692), .A2(n3115), .B1(n3116), .B2(n3092), .ZN(
        p8_muxs_out_2__17_) );
  AOI21_X1 U3323 ( .B1(reg3_reg[4]), .B2(reg3_reg[3]), .A(
        p8_minus_A_shifted_38_), .ZN(n3117) );
  OAI21_X1 U3324 ( .B1(reg3_reg[4]), .B2(reg3_reg[3]), .A(n2853), .ZN(n3118)
         );
  OAI22_X1 U3325 ( .A1(n3117), .A2(n2853), .B1(p8_minus_A_shifted_38_), .B2(
        n3118), .ZN(p8_muxs_out_2__18_) );
  NAND2_X1 U3326 ( .A1(B2[0]), .A2(n3120), .ZN(n3121) );
  XNOR2_X1 U3327 ( .A(n3121), .B(p8_Partial_products_sum_add_23_B_0_), .ZN(
        p8_muxs_out_3__6_) );
  OAI221_X1 U3328 ( .B1(B2[0]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_13_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3122) );
  OAI221_X1 U3329 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[1]), .C1(
        n2800), .C2(p8_minus_A_shifted_14_), .A(n3120), .ZN(n3123) );
  NAND2_X1 U3330 ( .A1(n3122), .A2(n3123), .ZN(p8_muxs_out_3__7_) );
  OAI221_X1 U3331 ( .B1(B2[1]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_14_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3124) );
  OAI221_X1 U3332 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[2]), .C1(
        n2800), .C2(p8_minus_A_shifted_15_), .A(n3120), .ZN(n3125) );
  NAND2_X1 U3333 ( .A1(n3124), .A2(n3125), .ZN(p8_muxs_out_3__8_) );
  OAI221_X1 U3334 ( .B1(B2[2]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_15_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3126) );
  OAI221_X1 U3335 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[3]), .C1(
        n2800), .C2(p8_minus_A_shifted_16_), .A(n3120), .ZN(n3127) );
  NAND2_X1 U3336 ( .A1(n3126), .A2(n3127), .ZN(p8_muxs_out_3__9_) );
  OAI221_X1 U3337 ( .B1(B2[3]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_16_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3128) );
  OAI221_X1 U3338 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[4]), .C1(
        n2800), .C2(p8_minus_A_shifted_17_), .A(n3120), .ZN(n3129) );
  NAND2_X1 U3339 ( .A1(n3128), .A2(n3129), .ZN(p8_muxs_out_3__10_) );
  OAI221_X1 U3340 ( .B1(B2[4]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_17_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3130) );
  OAI221_X1 U3341 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[5]), .C1(
        n2800), .C2(p8_minus_A_shifted_18_), .A(n3120), .ZN(n3131) );
  NAND2_X1 U3342 ( .A1(n3130), .A2(n3131), .ZN(p8_muxs_out_3__11_) );
  OAI221_X1 U3343 ( .B1(B2[5]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_18_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3132) );
  OAI221_X1 U3344 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[6]), .C1(
        n2800), .C2(p8_minus_A_shifted_19_), .A(n3120), .ZN(n3133) );
  NAND2_X1 U3345 ( .A1(n3132), .A2(n3133), .ZN(p8_muxs_out_3__12_) );
  OAI221_X1 U3346 ( .B1(B2[6]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_19_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3134) );
  OAI221_X1 U3347 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[7]), .C1(
        n2800), .C2(p8_minus_A_shifted_20_), .A(n3120), .ZN(n3135) );
  NAND2_X1 U3348 ( .A1(n3134), .A2(n3135), .ZN(p8_muxs_out_3__13_) );
  OAI221_X1 U3349 ( .B1(B2[7]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_20_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3136) );
  OAI221_X1 U3350 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[8]), .C1(
        n2800), .C2(p8_minus_A_shifted_21_), .A(n3120), .ZN(n3137) );
  NAND2_X1 U3351 ( .A1(n3136), .A2(n3137), .ZN(p8_muxs_out_3__14_) );
  OAI221_X1 U3352 ( .B1(B2[8]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_21_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3138) );
  OAI221_X1 U3353 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[9]), .C1(
        n2800), .C2(p8_minus_A_shifted_22_), .A(n3120), .ZN(n3139) );
  NAND2_X1 U3354 ( .A1(n3138), .A2(n3139), .ZN(p8_muxs_out_3__15_) );
  OAI221_X1 U3355 ( .B1(B2[9]), .B2(p8_Partial_products_sum_add_23_B_0_), .C1(
        p8_minus_A_shifted_22_), .C2(reg3_reg[6]), .A(n3119), .ZN(n3140) );
  OAI221_X1 U3356 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[10]), 
        .C1(n2800), .C2(p8_minus_A_shifted_23_), .A(n3120), .ZN(n3141) );
  NAND2_X1 U3357 ( .A1(n3140), .A2(n3141), .ZN(p8_muxs_out_3__16_) );
  OAI221_X1 U3358 ( .B1(B2[10]), .B2(p8_Partial_products_sum_add_23_B_0_), 
        .C1(p8_minus_A_shifted_23_), .C2(reg3_reg[6]), .A(n2686), .ZN(n3142)
         );
  OAI221_X1 U3359 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[11]), 
        .C1(n2800), .C2(n3068), .A(n3120), .ZN(n3143) );
  NAND2_X1 U3360 ( .A1(n3142), .A2(n3143), .ZN(p8_muxs_out_3__17_) );
  OAI221_X1 U3361 ( .B1(B2[11]), .B2(p8_Partial_products_sum_add_23_B_0_), 
        .C1(n3068), .C2(reg3_reg[6]), .A(n2686), .ZN(n3144) );
  OAI221_X1 U3362 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[12]), 
        .C1(n2800), .C2(p8_minus_A_shifted_25_), .A(n3120), .ZN(n3145) );
  NAND2_X1 U3363 ( .A1(n3144), .A2(n3145), .ZN(p8_muxs_out_3__18_) );
  OAI221_X1 U3364 ( .B1(B2[12]), .B2(p8_Partial_products_sum_add_23_B_0_), 
        .C1(p8_minus_A_shifted_25_), .C2(reg3_reg[6]), .A(n2686), .ZN(n3146)
         );
  OAI221_X1 U3365 ( .B1(p8_Partial_products_sum_add_23_B_0_), .B2(B2[13]), 
        .C1(n2800), .C2(p8_minus_A_shifted_38_), .A(n3120), .ZN(n3147) );
  NAND2_X1 U3366 ( .A1(n3146), .A2(n3147), .ZN(p8_muxs_out_3__19_) );
  AOI21_X1 U3367 ( .B1(reg3_reg[6]), .B2(reg3_reg[5]), .A(
        p8_minus_A_shifted_38_), .ZN(n3148) );
  OAI21_X1 U3368 ( .B1(reg3_reg[6]), .B2(reg3_reg[5]), .A(n2800), .ZN(n3149)
         );
  OAI22_X1 U3369 ( .A1(n3148), .A2(n2800), .B1(p8_minus_A_shifted_38_), .B2(
        n3149), .ZN(p8_muxs_out_3__20_) );
  AOI22_X1 U3370 ( .A1(reg4_reg[2]), .A2(reg4_reg[1]), .B1(n2841), .B2(n2795), 
        .ZN(n3150) );
  OAI221_X1 U3371 ( .B1(p9_minus_A_shifted_16_), .B2(reg4_reg[2]), .C1(B3[3]), 
        .C2(reg4_reg[3]), .A(n3151), .ZN(n3153) );
  OAI221_X1 U3372 ( .B1(reg4_reg[3]), .B2(B3[4]), .C1(n2847), .C2(
        p9_minus_A_shifted_17_), .A(n3150), .ZN(n3154) );
  NAND2_X1 U3373 ( .A1(n3153), .A2(n3154), .ZN(p9_muxs_out_1__6_) );
  OAI221_X1 U3374 ( .B1(B3[4]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_17_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3155) );
  OAI221_X1 U3375 ( .B1(reg4_reg[3]), .B2(B3[5]), .C1(n2847), .C2(
        p9_minus_A_shifted_18_), .A(n3150), .ZN(n3156) );
  OAI221_X1 U3376 ( .B1(B3[5]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_18_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3157) );
  OAI221_X1 U3377 ( .B1(reg4_reg[3]), .B2(B3[6]), .C1(n2847), .C2(
        p9_minus_A_shifted_19_), .A(n3150), .ZN(n3158) );
  NAND2_X1 U3378 ( .A1(n3157), .A2(n3158), .ZN(p9_muxs_out_1__8_) );
  OAI221_X1 U3379 ( .B1(B3[6]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_19_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3159) );
  OAI221_X1 U3380 ( .B1(reg4_reg[3]), .B2(B3[7]), .C1(n2847), .C2(
        p9_minus_A_shifted_20_), .A(n3150), .ZN(n3160) );
  NAND2_X1 U3381 ( .A1(n3159), .A2(n3160), .ZN(p9_muxs_out_1__9_) );
  OAI221_X1 U3382 ( .B1(B3[7]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_20_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3161) );
  OAI221_X1 U3383 ( .B1(reg4_reg[3]), .B2(B3[8]), .C1(n2847), .C2(
        p9_minus_A_shifted_21_), .A(n3150), .ZN(n3162) );
  NAND2_X1 U3384 ( .A1(n3161), .A2(n3162), .ZN(p9_muxs_out_1__10_) );
  OAI221_X1 U3385 ( .B1(B3[8]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_21_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3163) );
  OAI221_X1 U3386 ( .B1(reg4_reg[3]), .B2(B3[9]), .C1(n2847), .C2(
        p9_minus_A_shifted_22_), .A(n3150), .ZN(n3164) );
  NAND2_X1 U3387 ( .A1(n3163), .A2(n3164), .ZN(p9_muxs_out_1__11_) );
  OAI221_X1 U3388 ( .B1(B3[9]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_22_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3165) );
  OAI221_X1 U3389 ( .B1(reg4_reg[3]), .B2(B3[10]), .C1(n2847), .C2(
        p9_minus_A_shifted_23_), .A(n3150), .ZN(n3166) );
  NAND2_X1 U3390 ( .A1(n3165), .A2(n3166), .ZN(p9_muxs_out_1__12_) );
  OAI221_X1 U3391 ( .B1(B3[10]), .B2(reg4_reg[3]), .C1(p9_minus_A_shifted_23_), 
        .C2(reg4_reg[2]), .A(n3151), .ZN(n3167) );
  OAI221_X1 U3392 ( .B1(reg4_reg[3]), .B2(B3[11]), .C1(n2847), .C2(n3152), .A(
        n3150), .ZN(n3168) );
  NAND2_X1 U3393 ( .A1(n3167), .A2(n3168), .ZN(p9_muxs_out_1__13_) );
  OAI221_X1 U3394 ( .B1(B3[11]), .B2(reg4_reg[3]), .C1(n3152), .C2(reg4_reg[2]), .A(n3151), .ZN(n3169) );
  OAI221_X1 U3395 ( .B1(reg4_reg[3]), .B2(B3[12]), .C1(n2847), .C2(
        p9_minus_A_shifted_25_), .A(n3150), .ZN(n3170) );
  NAND2_X1 U3396 ( .A1(n3169), .A2(n3170), .ZN(p9_muxs_out_1__14_) );
  AOI22_X1 U3397 ( .A1(reg4_reg[3]), .A2(p9_minus_A_shifted_38_), .B1(B3[13]), 
        .B2(n2847), .ZN(n3171) );
  AOI22_X1 U3398 ( .A1(B3[12]), .A2(reg4_reg[2]), .B1(reg4_reg[3]), .B2(
        p9_minus_A_shifted_25_), .ZN(n3172) );
  AOI22_X1 U3399 ( .A1(n3150), .A2(n3171), .B1(n3172), .B2(n3151), .ZN(
        p9_muxs_out_1__15_) );
  AOI21_X1 U3400 ( .B1(reg4_reg[2]), .B2(reg4_reg[1]), .A(
        p9_minus_A_shifted_38_), .ZN(n3173) );
  OAI21_X1 U3401 ( .B1(reg4_reg[2]), .B2(reg4_reg[1]), .A(n2847), .ZN(n3174)
         );
  OAI22_X1 U3402 ( .A1(n3173), .A2(n2847), .B1(p9_minus_A_shifted_38_), .B2(
        n3174), .ZN(p9_muxs_out_1__16_) );
  AOI22_X1 U3403 ( .A1(reg4_reg[4]), .A2(reg4_reg[3]), .B1(n2847), .B2(n2829), 
        .ZN(n3175) );
  OAI221_X1 U3404 ( .B1(p9_minus_A_shifted_14_), .B2(reg4_reg[4]), .C1(B3[1]), 
        .C2(reg4_reg[5]), .A(n3176), .ZN(n3177) );
  OAI221_X1 U3405 ( .B1(reg4_reg[5]), .B2(B3[2]), .C1(n2854), .C2(
        p9_minus_A_shifted_15_), .A(n3175), .ZN(n3178) );
  NAND2_X1 U3406 ( .A1(n3177), .A2(n3178), .ZN(p9_muxs_out_2__6_) );
  OAI221_X1 U3407 ( .B1(B3[2]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_15_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3179) );
  OAI221_X1 U3408 ( .B1(reg4_reg[5]), .B2(B3[3]), .C1(n2854), .C2(
        p9_minus_A_shifted_16_), .A(n3175), .ZN(n3180) );
  NAND2_X1 U3409 ( .A1(n3179), .A2(n3180), .ZN(p9_muxs_out_2__7_) );
  OAI221_X1 U3410 ( .B1(B3[3]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_16_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3181) );
  OAI221_X1 U3411 ( .B1(reg4_reg[5]), .B2(B3[4]), .C1(n2854), .C2(
        p9_minus_A_shifted_17_), .A(n3175), .ZN(n3182) );
  NAND2_X1 U3412 ( .A1(n3181), .A2(n3182), .ZN(p9_muxs_out_2__8_) );
  OAI221_X1 U3413 ( .B1(B3[4]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_17_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3183) );
  OAI221_X1 U3414 ( .B1(reg4_reg[5]), .B2(B3[5]), .C1(n2854), .C2(
        p9_minus_A_shifted_18_), .A(n3175), .ZN(n3184) );
  NAND2_X1 U3415 ( .A1(n3183), .A2(n3184), .ZN(p9_muxs_out_2__9_) );
  OAI221_X1 U3416 ( .B1(B3[5]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_18_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3185) );
  OAI221_X1 U3417 ( .B1(reg4_reg[5]), .B2(B3[6]), .C1(n2854), .C2(
        p9_minus_A_shifted_19_), .A(n3175), .ZN(n3186) );
  NAND2_X1 U3418 ( .A1(n3185), .A2(n3186), .ZN(p9_muxs_out_2__10_) );
  OAI221_X1 U3419 ( .B1(B3[6]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_19_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3187) );
  OAI221_X1 U3420 ( .B1(reg4_reg[5]), .B2(B3[7]), .C1(n2854), .C2(
        p9_minus_A_shifted_20_), .A(n3175), .ZN(n3188) );
  NAND2_X1 U3421 ( .A1(n3187), .A2(n3188), .ZN(p9_muxs_out_2__11_) );
  OAI221_X1 U3422 ( .B1(B3[7]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_20_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3189) );
  OAI221_X1 U3423 ( .B1(reg4_reg[5]), .B2(B3[8]), .C1(n2854), .C2(
        p9_minus_A_shifted_21_), .A(n3175), .ZN(n3190) );
  NAND2_X1 U3424 ( .A1(n3189), .A2(n3190), .ZN(p9_muxs_out_2__12_) );
  OAI221_X1 U3425 ( .B1(B3[8]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_21_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3191) );
  OAI221_X1 U3426 ( .B1(reg4_reg[5]), .B2(B3[9]), .C1(n2854), .C2(
        p9_minus_A_shifted_22_), .A(n3175), .ZN(n3192) );
  NAND2_X1 U3427 ( .A1(n3191), .A2(n3192), .ZN(p9_muxs_out_2__13_) );
  OAI221_X1 U3428 ( .B1(B3[9]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_22_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3193) );
  OAI221_X1 U3429 ( .B1(reg4_reg[5]), .B2(B3[10]), .C1(n2854), .C2(
        p9_minus_A_shifted_23_), .A(n3175), .ZN(n3194) );
  NAND2_X1 U3430 ( .A1(n3193), .A2(n3194), .ZN(p9_muxs_out_2__14_) );
  OAI221_X1 U3431 ( .B1(B3[10]), .B2(reg4_reg[5]), .C1(p9_minus_A_shifted_23_), 
        .C2(reg4_reg[4]), .A(n3176), .ZN(n3195) );
  OAI221_X1 U3432 ( .B1(reg4_reg[5]), .B2(B3[11]), .C1(n2854), .C2(n3152), .A(
        n3175), .ZN(n3196) );
  NAND2_X1 U3433 ( .A1(n3195), .A2(n3196), .ZN(p9_muxs_out_2__15_) );
  OAI221_X1 U3434 ( .B1(B3[11]), .B2(reg4_reg[5]), .C1(n3152), .C2(reg4_reg[4]), .A(n3176), .ZN(n3197) );
  OAI221_X1 U3435 ( .B1(reg4_reg[5]), .B2(B3[12]), .C1(n2854), .C2(
        p9_minus_A_shifted_25_), .A(n2693), .ZN(n3198) );
  NAND2_X1 U3436 ( .A1(n3197), .A2(n3198), .ZN(p9_muxs_out_2__16_) );
  AOI22_X1 U3437 ( .A1(reg4_reg[5]), .A2(p9_minus_A_shifted_38_), .B1(B3[13]), 
        .B2(n2854), .ZN(n3199) );
  AOI22_X1 U3438 ( .A1(B3[12]), .A2(reg4_reg[4]), .B1(reg4_reg[5]), .B2(
        p9_minus_A_shifted_25_), .ZN(n3200) );
  AOI22_X1 U3439 ( .A1(n2693), .A2(n3199), .B1(n3200), .B2(n3176), .ZN(
        p9_muxs_out_2__17_) );
  AOI21_X1 U3440 ( .B1(reg4_reg[4]), .B2(reg4_reg[3]), .A(
        p9_minus_A_shifted_38_), .ZN(n3201) );
  OAI21_X1 U3441 ( .B1(reg4_reg[4]), .B2(reg4_reg[3]), .A(n2854), .ZN(n3202)
         );
  OAI22_X1 U3442 ( .A1(n3201), .A2(n2854), .B1(p9_minus_A_shifted_38_), .B2(
        n3202), .ZN(p9_muxs_out_2__18_) );
  NAND2_X1 U3443 ( .A1(B3[0]), .A2(n3204), .ZN(n3205) );
  XNOR2_X1 U3444 ( .A(n3205), .B(p9_Partial_products_sum_add_23_B_0_), .ZN(
        p9_muxs_out_3__6_) );
  OAI221_X1 U3445 ( .B1(B3[0]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_13_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3206) );
  OAI221_X1 U3446 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[1]), .C1(
        n2801), .C2(p9_minus_A_shifted_14_), .A(n3204), .ZN(n3207) );
  NAND2_X1 U3447 ( .A1(n3206), .A2(n3207), .ZN(p9_muxs_out_3__7_) );
  OAI221_X1 U3448 ( .B1(B3[1]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_14_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3208) );
  OAI221_X1 U3449 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[2]), .C1(
        n2801), .C2(p9_minus_A_shifted_15_), .A(n3204), .ZN(n3209) );
  NAND2_X1 U3450 ( .A1(n3208), .A2(n3209), .ZN(p9_muxs_out_3__8_) );
  OAI221_X1 U3451 ( .B1(B3[2]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_15_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3210) );
  OAI221_X1 U3452 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[3]), .C1(
        n2801), .C2(p9_minus_A_shifted_16_), .A(n3204), .ZN(n3211) );
  NAND2_X1 U3453 ( .A1(n3210), .A2(n3211), .ZN(p9_muxs_out_3__9_) );
  OAI221_X1 U3454 ( .B1(B3[3]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_16_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3212) );
  OAI221_X1 U3455 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[4]), .C1(
        n2801), .C2(p9_minus_A_shifted_17_), .A(n3204), .ZN(n3213) );
  NAND2_X1 U3456 ( .A1(n3212), .A2(n3213), .ZN(p9_muxs_out_3__10_) );
  OAI221_X1 U3457 ( .B1(B3[4]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_17_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3214) );
  OAI221_X1 U3458 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[5]), .C1(
        n2801), .C2(p9_minus_A_shifted_18_), .A(n3204), .ZN(n3215) );
  NAND2_X1 U3459 ( .A1(n3214), .A2(n3215), .ZN(p9_muxs_out_3__11_) );
  OAI221_X1 U3460 ( .B1(B3[5]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_18_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3216) );
  OAI221_X1 U3461 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[6]), .C1(
        n2801), .C2(p9_minus_A_shifted_19_), .A(n3204), .ZN(n3217) );
  NAND2_X1 U3462 ( .A1(n3216), .A2(n3217), .ZN(p9_muxs_out_3__12_) );
  OAI221_X1 U3463 ( .B1(B3[6]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_19_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3218) );
  OAI221_X1 U3464 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[7]), .C1(
        n2801), .C2(p9_minus_A_shifted_20_), .A(n3204), .ZN(n3219) );
  NAND2_X1 U3465 ( .A1(n3218), .A2(n3219), .ZN(p9_muxs_out_3__13_) );
  OAI221_X1 U3466 ( .B1(B3[7]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_20_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3220) );
  OAI221_X1 U3467 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[8]), .C1(
        n2801), .C2(p9_minus_A_shifted_21_), .A(n3204), .ZN(n3221) );
  NAND2_X1 U3468 ( .A1(n3220), .A2(n3221), .ZN(p9_muxs_out_3__14_) );
  OAI221_X1 U3469 ( .B1(B3[8]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_21_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3222) );
  OAI221_X1 U3470 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[9]), .C1(
        n2801), .C2(p9_minus_A_shifted_22_), .A(n3204), .ZN(n3223) );
  NAND2_X1 U3471 ( .A1(n3222), .A2(n3223), .ZN(p9_muxs_out_3__15_) );
  OAI221_X1 U3472 ( .B1(B3[9]), .B2(p9_Partial_products_sum_add_23_B_0_), .C1(
        p9_minus_A_shifted_22_), .C2(reg4_reg[6]), .A(n3203), .ZN(n3224) );
  OAI221_X1 U3473 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[10]), 
        .C1(n2801), .C2(p9_minus_A_shifted_23_), .A(n3204), .ZN(n3225) );
  NAND2_X1 U3474 ( .A1(n3224), .A2(n3225), .ZN(p9_muxs_out_3__16_) );
  OAI221_X1 U3475 ( .B1(B3[10]), .B2(p9_Partial_products_sum_add_23_B_0_), 
        .C1(p9_minus_A_shifted_23_), .C2(reg4_reg[6]), .A(n2688), .ZN(n3226)
         );
  OAI221_X1 U3476 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[11]), 
        .C1(n2801), .C2(n3152), .A(n3204), .ZN(n3227) );
  NAND2_X1 U3477 ( .A1(n3226), .A2(n3227), .ZN(p9_muxs_out_3__17_) );
  OAI221_X1 U3478 ( .B1(B3[11]), .B2(p9_Partial_products_sum_add_23_B_0_), 
        .C1(n3152), .C2(reg4_reg[6]), .A(n2688), .ZN(n3228) );
  OAI221_X1 U3479 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[12]), 
        .C1(n2801), .C2(p9_minus_A_shifted_25_), .A(n3204), .ZN(n3229) );
  NAND2_X1 U3480 ( .A1(n3228), .A2(n3229), .ZN(p9_muxs_out_3__18_) );
  OAI221_X1 U3481 ( .B1(B3[12]), .B2(p9_Partial_products_sum_add_23_B_0_), 
        .C1(p9_minus_A_shifted_25_), .C2(reg4_reg[6]), .A(n2688), .ZN(n3230)
         );
  OAI221_X1 U3482 ( .B1(p9_Partial_products_sum_add_23_B_0_), .B2(B3[13]), 
        .C1(n2801), .C2(p9_minus_A_shifted_38_), .A(n3204), .ZN(n3231) );
  NAND2_X1 U3483 ( .A1(n3230), .A2(n3231), .ZN(p9_muxs_out_3__19_) );
  AOI21_X1 U3484 ( .B1(reg4_reg[6]), .B2(reg4_reg[5]), .A(
        p9_minus_A_shifted_38_), .ZN(n3232) );
  OAI21_X1 U3485 ( .B1(reg4_reg[6]), .B2(reg4_reg[5]), .A(n2801), .ZN(n3233)
         );
  OAI22_X1 U3486 ( .A1(n3232), .A2(n2801), .B1(p9_minus_A_shifted_38_), .B2(
        n3233), .ZN(p9_muxs_out_3__20_) );
  OAI221_X1 U3487 ( .B1(p11_minus_A_shifted_16_), .B2(A1[2]), .C1(reg2[3]), 
        .C2(A1[3]), .A(n3235), .ZN(n3236) );
  OAI221_X1 U3488 ( .B1(A1[3]), .B2(reg2[4]), .C1(n3259), .C2(n2817), .A(n3260), .ZN(n3237) );
  NAND2_X1 U3489 ( .A1(n3236), .A2(n3237), .ZN(p11_muxs_out_1__6_) );
  OAI221_X1 U3490 ( .B1(reg2[4]), .B2(A1[3]), .C1(n2817), .C2(A1[2]), .A(n3235), .ZN(n3238) );
  OAI221_X1 U3491 ( .B1(A1[3]), .B2(reg2[5]), .C1(n3258), .C2(n2834), .A(n3260), .ZN(n3239) );
  OAI221_X1 U3492 ( .B1(reg2[5]), .B2(A1[3]), .C1(n2834), .C2(A1[2]), .A(n3235), .ZN(n3240) );
  OAI221_X1 U3493 ( .B1(A1[3]), .B2(reg2[6]), .C1(n3258), .C2(n2835), .A(n3260), .ZN(n3241) );
  NAND2_X1 U3494 ( .A1(n3240), .A2(n3241), .ZN(p11_muxs_out_1__8_) );
  OAI221_X1 U3495 ( .B1(reg2[6]), .B2(A1[3]), .C1(n2835), .C2(A1[2]), .A(n3235), .ZN(n3242) );
  OAI221_X1 U3496 ( .B1(A1[3]), .B2(reg2[7]), .C1(n3258), .C2(n2831), .A(n3260), .ZN(n3243) );
  NAND2_X1 U3497 ( .A1(n3242), .A2(n3243), .ZN(p11_muxs_out_1__9_) );
  OAI221_X1 U3498 ( .B1(reg2[7]), .B2(A1[3]), .C1(n2831), .C2(A1[2]), .A(n3235), .ZN(n3244) );
  OAI221_X1 U3499 ( .B1(A1[3]), .B2(reg2[8]), .C1(n3259), .C2(n2811), .A(n3260), .ZN(n3245) );
  NAND2_X1 U3500 ( .A1(n3244), .A2(n3245), .ZN(p11_muxs_out_1__10_) );
  OAI221_X1 U3501 ( .B1(reg2[8]), .B2(A1[3]), .C1(n2811), .C2(A1[2]), .A(n3235), .ZN(n3246) );
  OAI221_X1 U3502 ( .B1(A1[3]), .B2(reg2[9]), .C1(n3259), .C2(n2816), .A(n3260), .ZN(n3247) );
  NAND2_X1 U3503 ( .A1(n3246), .A2(n3247), .ZN(p11_muxs_out_1__11_) );
  OAI221_X1 U3504 ( .B1(reg2[9]), .B2(A1[3]), .C1(n2816), .C2(A1[2]), .A(n3235), .ZN(n3248) );
  OAI221_X1 U3505 ( .B1(A1[3]), .B2(reg2[10]), .C1(n3259), .C2(n2833), .A(
        n3260), .ZN(n3249) );
  NAND2_X1 U3506 ( .A1(n3248), .A2(n3249), .ZN(p11_muxs_out_1__12_) );
  OAI221_X1 U3507 ( .B1(reg2[10]), .B2(A1[3]), .C1(n2833), .C2(A1[2]), .A(
        n3235), .ZN(n3250) );
  OAI221_X1 U3508 ( .B1(A1[3]), .B2(reg2[11]), .C1(n3259), .C2(n2862), .A(
        n3260), .ZN(n3251) );
  NAND2_X1 U3509 ( .A1(n3250), .A2(n3251), .ZN(p11_muxs_out_1__13_) );
  OAI221_X1 U3510 ( .B1(reg2[11]), .B2(A1[3]), .C1(n2862), .C2(A1[2]), .A(
        n3235), .ZN(n3252) );
  OAI221_X1 U3511 ( .B1(A1[3]), .B2(reg2[12]), .C1(n3259), .C2(n2863), .A(
        n3260), .ZN(n3253) );
  NAND2_X1 U3512 ( .A1(n3252), .A2(n3253), .ZN(p11_muxs_out_1__14_) );
  AOI22_X1 U3513 ( .A1(A1[3]), .A2(n2860), .B1(reg2[13]), .B2(n3259), .ZN(
        n3254) );
  AOI22_X1 U3514 ( .A1(reg2[12]), .A2(A1[2]), .B1(A1[3]), .B2(n2863), .ZN(
        n3255) );
  AOI22_X1 U3515 ( .A1(n3260), .A2(n3254), .B1(n3255), .B2(n3235), .ZN(
        p11_muxs_out_1__15_) );
  AOI21_X1 U3516 ( .B1(A1[2]), .B2(A1[1]), .A(n2860), .ZN(n3256) );
  OAI21_X1 U3517 ( .B1(A1[2]), .B2(A1[1]), .A(n3259), .ZN(n3257) );
  OAI22_X1 U3518 ( .A1(n3256), .A2(n3259), .B1(n2860), .B2(n3257), .ZN(
        p11_muxs_out_1__16_) );
  OAI221_X1 U3519 ( .B1(p11_minus_A_shifted_14_), .B2(A1[4]), .C1(reg2[1]), 
        .C2(A1[5]), .A(n3263), .ZN(n3264) );
  OAI221_X1 U3520 ( .B1(A1[5]), .B2(reg2[2]), .C1(n3290), .C2(n2820), .A(n3262), .ZN(n3265) );
  NAND2_X1 U3521 ( .A1(n3264), .A2(n3265), .ZN(p11_muxs_out_2__6_) );
  OAI221_X1 U3522 ( .B1(reg2[2]), .B2(A1[5]), .C1(n2820), .C2(A1[4]), .A(n3263), .ZN(n3266) );
  OAI221_X1 U3523 ( .B1(A1[5]), .B2(reg2[3]), .C1(n3290), .C2(
        p11_minus_A_shifted_16_), .A(n3262), .ZN(n3267) );
  NAND2_X1 U3524 ( .A1(n3266), .A2(n3267), .ZN(p11_muxs_out_2__7_) );
  OAI221_X1 U3525 ( .B1(reg2[3]), .B2(A1[5]), .C1(p11_minus_A_shifted_16_), 
        .C2(A1[4]), .A(n3263), .ZN(n3268) );
  OAI221_X1 U3526 ( .B1(A1[5]), .B2(reg2[4]), .C1(n3290), .C2(n2817), .A(n3262), .ZN(n3269) );
  OAI221_X1 U3527 ( .B1(reg2[4]), .B2(A1[5]), .C1(n2817), .C2(A1[4]), .A(n3263), .ZN(n3270) );
  OAI221_X1 U3528 ( .B1(A1[5]), .B2(reg2[5]), .C1(n3290), .C2(n2834), .A(n3262), .ZN(n3271) );
  NAND2_X1 U3529 ( .A1(n3270), .A2(n3271), .ZN(p11_muxs_out_2__9_) );
  OAI221_X1 U3530 ( .B1(reg2[5]), .B2(A1[5]), .C1(n2834), .C2(A1[4]), .A(n3263), .ZN(n3272) );
  OAI221_X1 U3531 ( .B1(A1[5]), .B2(reg2[6]), .C1(n3290), .C2(n2835), .A(n3262), .ZN(n3273) );
  NAND2_X1 U3532 ( .A1(n3272), .A2(n3273), .ZN(p11_muxs_out_2__10_) );
  OAI221_X1 U3533 ( .B1(reg2[6]), .B2(A1[5]), .C1(n2835), .C2(A1[4]), .A(n3263), .ZN(n3274) );
  OAI221_X1 U3534 ( .B1(A1[5]), .B2(reg2[7]), .C1(n3290), .C2(n2831), .A(n3262), .ZN(n3275) );
  NAND2_X1 U3535 ( .A1(n3274), .A2(n3275), .ZN(p11_muxs_out_2__11_) );
  OAI221_X1 U3536 ( .B1(reg2[7]), .B2(A1[5]), .C1(n2831), .C2(A1[4]), .A(n3263), .ZN(n3276) );
  OAI221_X1 U3537 ( .B1(A1[5]), .B2(reg2[8]), .C1(n3290), .C2(n2811), .A(n3262), .ZN(n3277) );
  NAND2_X1 U3538 ( .A1(n3276), .A2(n3277), .ZN(p11_muxs_out_2__12_) );
  OAI221_X1 U3539 ( .B1(reg2[8]), .B2(A1[5]), .C1(n2811), .C2(A1[4]), .A(n3263), .ZN(n3278) );
  OAI221_X1 U3540 ( .B1(A1[5]), .B2(reg2[9]), .C1(n3290), .C2(n2816), .A(n3262), .ZN(n3279) );
  NAND2_X1 U3541 ( .A1(n3278), .A2(n3279), .ZN(p11_muxs_out_2__13_) );
  OAI221_X1 U3542 ( .B1(reg2[9]), .B2(A1[5]), .C1(n2816), .C2(A1[4]), .A(n3263), .ZN(n3280) );
  OAI221_X1 U3543 ( .B1(A1[5]), .B2(reg2[10]), .C1(n3290), .C2(n2833), .A(
        n3262), .ZN(n3281) );
  NAND2_X1 U3544 ( .A1(n3280), .A2(n3281), .ZN(p11_muxs_out_2__14_) );
  OAI221_X1 U3545 ( .B1(reg2[10]), .B2(A1[5]), .C1(n2833), .C2(A1[4]), .A(
        n3263), .ZN(n3282) );
  OAI221_X1 U3546 ( .B1(A1[5]), .B2(reg2[11]), .C1(n3290), .C2(n2862), .A(
        n3262), .ZN(n3283) );
  NAND2_X1 U3547 ( .A1(n3282), .A2(n3283), .ZN(p11_muxs_out_2__15_) );
  OAI221_X1 U3548 ( .B1(reg2[11]), .B2(A1[5]), .C1(n2862), .C2(A1[4]), .A(
        n3263), .ZN(n3284) );
  OAI221_X1 U3549 ( .B1(A1[5]), .B2(reg2[12]), .C1(n3290), .C2(n2863), .A(
        n3262), .ZN(n3285) );
  NAND2_X1 U3550 ( .A1(n3284), .A2(n3285), .ZN(p11_muxs_out_2__16_) );
  AOI22_X1 U3551 ( .A1(A1[5]), .A2(n2860), .B1(reg2[13]), .B2(n3290), .ZN(
        n3286) );
  AOI22_X1 U3552 ( .A1(reg2[12]), .A2(A1[4]), .B1(A1[5]), .B2(n2863), .ZN(
        n3287) );
  AOI22_X1 U3553 ( .A1(n3262), .A2(n3286), .B1(n3287), .B2(n3263), .ZN(
        p11_muxs_out_2__17_) );
  AOI21_X1 U3554 ( .B1(A1[4]), .B2(A1[3]), .A(n2860), .ZN(n3288) );
  OAI21_X1 U3555 ( .B1(A1[4]), .B2(A1[3]), .A(n3290), .ZN(n3289) );
  OAI22_X1 U3556 ( .A1(n3288), .A2(n3290), .B1(n2860), .B2(n3289), .ZN(
        p11_muxs_out_2__18_) );
  NAND2_X1 U3557 ( .A1(reg2[0]), .A2(n3293), .ZN(n3294) );
  XNOR2_X1 U3558 ( .A(n3294), .B(n3324), .ZN(p11_muxs_out_3__6_) );
  OAI221_X1 U3559 ( .B1(reg2[0]), .B2(n3324), .C1(n2838), .C2(A1[6]), .A(n3292), .ZN(n3295) );
  OAI221_X1 U3560 ( .B1(n3324), .B2(reg2[1]), .C1(n3323), .C2(
        p11_minus_A_shifted_14_), .A(n3293), .ZN(n3296) );
  NAND2_X1 U3561 ( .A1(n3295), .A2(n3296), .ZN(p11_muxs_out_3__7_) );
  OAI221_X1 U3562 ( .B1(reg2[1]), .B2(n3324), .C1(p11_minus_A_shifted_14_), 
        .C2(A1[6]), .A(n3292), .ZN(n3297) );
  OAI221_X1 U3563 ( .B1(n3324), .B2(reg2[2]), .C1(n3323), .C2(n2820), .A(n3293), .ZN(n3298) );
  NAND2_X1 U3564 ( .A1(n3297), .A2(n3298), .ZN(p11_muxs_out_3__8_) );
  OAI221_X1 U3565 ( .B1(reg2[2]), .B2(n3324), .C1(n2820), .C2(A1[6]), .A(n3292), .ZN(n3299) );
  OAI221_X1 U3566 ( .B1(n3324), .B2(reg2[3]), .C1(n3323), .C2(
        p11_minus_A_shifted_16_), .A(n3293), .ZN(n3300) );
  NAND2_X1 U3567 ( .A1(n3299), .A2(n3300), .ZN(p11_muxs_out_3__9_) );
  OAI221_X1 U3568 ( .B1(reg2[3]), .B2(n3324), .C1(p11_minus_A_shifted_16_), 
        .C2(A1[6]), .A(n3292), .ZN(n3301) );
  OAI221_X1 U3569 ( .B1(n3324), .B2(reg2[4]), .C1(n3323), .C2(n2817), .A(n3293), .ZN(n3302) );
  NAND2_X1 U3570 ( .A1(n3301), .A2(n3302), .ZN(p11_muxs_out_3__10_) );
  OAI221_X1 U3571 ( .B1(reg2[4]), .B2(n3324), .C1(n2817), .C2(A1[6]), .A(n3292), .ZN(n3303) );
  OAI221_X1 U3572 ( .B1(n3324), .B2(reg2[5]), .C1(n3323), .C2(n2834), .A(n3293), .ZN(n3304) );
  NAND2_X1 U3573 ( .A1(n3303), .A2(n3304), .ZN(p11_muxs_out_3__11_) );
  OAI221_X1 U3574 ( .B1(reg2[5]), .B2(n3324), .C1(n2834), .C2(A1[6]), .A(n3292), .ZN(n3305) );
  OAI221_X1 U3575 ( .B1(n3324), .B2(reg2[6]), .C1(n3323), .C2(n2835), .A(n3293), .ZN(n3306) );
  NAND2_X1 U3576 ( .A1(n3305), .A2(n3306), .ZN(p11_muxs_out_3__12_) );
  OAI221_X1 U3577 ( .B1(reg2[6]), .B2(n3324), .C1(n2835), .C2(A1[6]), .A(n3292), .ZN(n3307) );
  OAI221_X1 U3578 ( .B1(n3324), .B2(reg2[7]), .C1(n3323), .C2(n2831), .A(n3293), .ZN(n3308) );
  NAND2_X1 U3579 ( .A1(n3307), .A2(n3308), .ZN(p11_muxs_out_3__13_) );
  OAI221_X1 U3580 ( .B1(reg2[7]), .B2(n3324), .C1(n2831), .C2(A1[6]), .A(n3292), .ZN(n3309) );
  OAI221_X1 U3581 ( .B1(n3324), .B2(reg2[8]), .C1(n3323), .C2(n2811), .A(n3293), .ZN(n3310) );
  NAND2_X1 U3582 ( .A1(n3309), .A2(n3310), .ZN(p11_muxs_out_3__14_) );
  OAI221_X1 U3583 ( .B1(reg2[8]), .B2(n3324), .C1(n2811), .C2(A1[6]), .A(n3292), .ZN(n3311) );
  OAI221_X1 U3584 ( .B1(n3324), .B2(reg2[9]), .C1(n3323), .C2(n2816), .A(n3293), .ZN(n3312) );
  NAND2_X1 U3585 ( .A1(n3311), .A2(n3312), .ZN(p11_muxs_out_3__15_) );
  OAI221_X1 U3586 ( .B1(reg2[9]), .B2(n3324), .C1(n2816), .C2(A1[6]), .A(n3326), .ZN(n3313) );
  OAI221_X1 U3587 ( .B1(n3324), .B2(reg2[10]), .C1(n3323), .C2(n2833), .A(
        n3293), .ZN(n3314) );
  NAND2_X1 U3588 ( .A1(n3313), .A2(n3314), .ZN(p11_muxs_out_3__16_) );
  OAI221_X1 U3589 ( .B1(reg2[10]), .B2(n3324), .C1(n2833), .C2(A1[6]), .A(
        n3326), .ZN(n3315) );
  OAI221_X1 U3590 ( .B1(n3324), .B2(reg2[11]), .C1(n3323), .C2(n2862), .A(
        n3293), .ZN(n3316) );
  NAND2_X1 U3591 ( .A1(n3315), .A2(n3316), .ZN(p11_muxs_out_3__17_) );
  OAI221_X1 U3592 ( .B1(reg2[11]), .B2(n3324), .C1(n2862), .C2(A1[6]), .A(
        n3326), .ZN(n3317) );
  OAI221_X1 U3593 ( .B1(n3324), .B2(reg2[12]), .C1(n3323), .C2(n2863), .A(
        n3293), .ZN(n3318) );
  NAND2_X1 U3594 ( .A1(n3317), .A2(n3318), .ZN(p11_muxs_out_3__18_) );
  OAI221_X1 U3595 ( .B1(reg2[12]), .B2(n3324), .C1(n2863), .C2(A1[6]), .A(
        n3326), .ZN(n3319) );
  OAI221_X1 U3596 ( .B1(n3324), .B2(reg2[13]), .C1(n3323), .C2(n2860), .A(
        n3293), .ZN(n3320) );
  AOI21_X1 U3597 ( .B1(A1[6]), .B2(A1[5]), .A(n2860), .ZN(n3321) );
  OAI21_X1 U3598 ( .B1(A1[6]), .B2(A1[5]), .A(n3323), .ZN(n3322) );
  OAI22_X1 U3599 ( .A1(n3321), .A2(n3323), .B1(n2860), .B2(n3322), .ZN(
        p11_muxs_out_3__20_) );
  OAI221_X1 U3600 ( .B1(p10_minus_A_shifted_16_), .B2(A2[2]), .C1(reg4[3]), 
        .C2(A2[3]), .A(n3330), .ZN(n3331) );
  OAI221_X1 U3601 ( .B1(A2[3]), .B2(reg4[4]), .C1(n3354), .C2(n2818), .A(n3329), .ZN(n3332) );
  NAND2_X1 U3602 ( .A1(n3331), .A2(n3332), .ZN(p10_muxs_out_1__6_) );
  OAI221_X1 U3603 ( .B1(reg4[4]), .B2(A2[3]), .C1(n2818), .C2(A2[2]), .A(n3330), .ZN(n3333) );
  OAI221_X1 U3604 ( .B1(A2[3]), .B2(reg4[5]), .C1(n3353), .C2(n2813), .A(n3329), .ZN(n3334) );
  OAI221_X1 U3605 ( .B1(reg4[5]), .B2(A2[3]), .C1(n2813), .C2(A2[2]), .A(n3330), .ZN(n3335) );
  OAI221_X1 U3606 ( .B1(A2[3]), .B2(reg4[6]), .C1(n3353), .C2(n2815), .A(n3355), .ZN(n3336) );
  NAND2_X1 U3607 ( .A1(n3335), .A2(n3336), .ZN(p10_muxs_out_1__8_) );
  OAI221_X1 U3608 ( .B1(reg4[6]), .B2(A2[3]), .C1(n2815), .C2(A2[2]), .A(n3330), .ZN(n3337) );
  OAI221_X1 U3609 ( .B1(A2[3]), .B2(reg4[7]), .C1(n3353), .C2(n2830), .A(n3355), .ZN(n3338) );
  NAND2_X1 U3610 ( .A1(n3337), .A2(n3338), .ZN(p10_muxs_out_1__9_) );
  OAI221_X1 U3611 ( .B1(reg4[7]), .B2(A2[3]), .C1(n2830), .C2(A2[2]), .A(n3330), .ZN(n3339) );
  OAI221_X1 U3612 ( .B1(A2[3]), .B2(reg4[8]), .C1(n3354), .C2(n2832), .A(n3329), .ZN(n3340) );
  NAND2_X1 U3613 ( .A1(n3339), .A2(n3340), .ZN(p10_muxs_out_1__10_) );
  OAI221_X1 U3614 ( .B1(reg4[8]), .B2(A2[3]), .C1(n2832), .C2(A2[2]), .A(n3330), .ZN(n3341) );
  OAI221_X1 U3615 ( .B1(A2[3]), .B2(reg4[9]), .C1(n3354), .C2(n2814), .A(n3355), .ZN(n3342) );
  NAND2_X1 U3616 ( .A1(n3341), .A2(n3342), .ZN(p10_muxs_out_1__11_) );
  OAI221_X1 U3617 ( .B1(reg4[9]), .B2(A2[3]), .C1(n2814), .C2(A2[2]), .A(n3330), .ZN(n3343) );
  OAI221_X1 U3618 ( .B1(A2[3]), .B2(reg4[10]), .C1(n3354), .C2(n2810), .A(
        n3355), .ZN(n3344) );
  NAND2_X1 U3619 ( .A1(n3343), .A2(n3344), .ZN(p10_muxs_out_1__12_) );
  OAI221_X1 U3620 ( .B1(reg4[10]), .B2(A2[3]), .C1(n2810), .C2(A2[2]), .A(
        n3330), .ZN(n3345) );
  OAI221_X1 U3621 ( .B1(A2[3]), .B2(reg4[11]), .C1(n3354), .C2(n2861), .A(
        n3355), .ZN(n3346) );
  NAND2_X1 U3622 ( .A1(n3345), .A2(n3346), .ZN(p10_muxs_out_1__13_) );
  OAI221_X1 U3623 ( .B1(reg4[11]), .B2(A2[3]), .C1(n2861), .C2(A2[2]), .A(
        n3330), .ZN(n3347) );
  OAI221_X1 U3624 ( .B1(A2[3]), .B2(reg4[12]), .C1(n3354), .C2(n2858), .A(
        n3355), .ZN(n3348) );
  NAND2_X1 U3625 ( .A1(n3347), .A2(n3348), .ZN(p10_muxs_out_1__14_) );
  AOI22_X1 U3626 ( .A1(A2[3]), .A2(n2859), .B1(reg4[13]), .B2(n3354), .ZN(
        n3349) );
  AOI22_X1 U3627 ( .A1(reg4[12]), .A2(A2[2]), .B1(A2[3]), .B2(n2858), .ZN(
        n3350) );
  AOI22_X1 U3628 ( .A1(n3355), .A2(n3349), .B1(n3350), .B2(n3330), .ZN(
        p10_muxs_out_1__15_) );
  AOI21_X1 U3629 ( .B1(A2[2]), .B2(A2[1]), .A(n2859), .ZN(n3351) );
  OAI21_X1 U3630 ( .B1(A2[2]), .B2(A2[1]), .A(n3354), .ZN(n3352) );
  OAI22_X1 U3631 ( .A1(n3351), .A2(n3354), .B1(n2859), .B2(n3352), .ZN(
        p10_muxs_out_1__16_) );
  OAI221_X1 U3632 ( .B1(p10_minus_A_shifted_14_), .B2(A2[4]), .C1(reg4[1]), 
        .C2(A2[5]), .A(n3384), .ZN(n3356) );
  OAI221_X1 U3633 ( .B1(A2[5]), .B2(reg4[2]), .C1(n3382), .C2(n2821), .A(n3383), .ZN(n3357) );
  NAND2_X1 U3634 ( .A1(n3356), .A2(n3357), .ZN(p10_muxs_out_2__6_) );
  OAI221_X1 U3635 ( .B1(reg4[2]), .B2(A2[5]), .C1(n2821), .C2(A2[4]), .A(n3384), .ZN(n3358) );
  OAI221_X1 U3636 ( .B1(A2[5]), .B2(reg4[3]), .C1(n3382), .C2(
        p10_minus_A_shifted_16_), .A(n3383), .ZN(n3359) );
  NAND2_X1 U3637 ( .A1(n3358), .A2(n3359), .ZN(p10_muxs_out_2__7_) );
  OAI221_X1 U3638 ( .B1(reg4[3]), .B2(A2[5]), .C1(p10_minus_A_shifted_16_), 
        .C2(A2[4]), .A(n3384), .ZN(n3360) );
  OAI221_X1 U3639 ( .B1(A2[5]), .B2(reg4[4]), .C1(n3382), .C2(n2818), .A(n3383), .ZN(n3361) );
  NAND2_X1 U3640 ( .A1(n3360), .A2(n3361), .ZN(p10_muxs_out_2__8_) );
  OAI221_X1 U3641 ( .B1(reg4[4]), .B2(A2[5]), .C1(n2818), .C2(A2[4]), .A(n3384), .ZN(n3362) );
  OAI221_X1 U3642 ( .B1(A2[5]), .B2(reg4[5]), .C1(n3382), .C2(n2813), .A(n3383), .ZN(n3363) );
  NAND2_X1 U3643 ( .A1(n3362), .A2(n3363), .ZN(p10_muxs_out_2__9_) );
  OAI221_X1 U3644 ( .B1(reg4[5]), .B2(A2[5]), .C1(n2813), .C2(A2[4]), .A(n3384), .ZN(n3364) );
  OAI221_X1 U3645 ( .B1(A2[5]), .B2(reg4[6]), .C1(n3382), .C2(n2815), .A(n3383), .ZN(n3365) );
  NAND2_X1 U3646 ( .A1(n3364), .A2(n3365), .ZN(p10_muxs_out_2__10_) );
  OAI221_X1 U3647 ( .B1(reg4[6]), .B2(A2[5]), .C1(n2815), .C2(A2[4]), .A(n3384), .ZN(n3366) );
  OAI221_X1 U3648 ( .B1(A2[5]), .B2(reg4[7]), .C1(n3382), .C2(n2830), .A(n3383), .ZN(n3367) );
  NAND2_X1 U3649 ( .A1(n3366), .A2(n3367), .ZN(p10_muxs_out_2__11_) );
  OAI221_X1 U3650 ( .B1(reg4[7]), .B2(A2[5]), .C1(n2830), .C2(A2[4]), .A(n3384), .ZN(n3368) );
  OAI221_X1 U3651 ( .B1(A2[5]), .B2(reg4[8]), .C1(n3382), .C2(n2832), .A(n3383), .ZN(n3369) );
  NAND2_X1 U3652 ( .A1(n3368), .A2(n3369), .ZN(p10_muxs_out_2__12_) );
  OAI221_X1 U3653 ( .B1(reg4[8]), .B2(A2[5]), .C1(n2832), .C2(A2[4]), .A(n3384), .ZN(n3370) );
  OAI221_X1 U3654 ( .B1(A2[5]), .B2(reg4[9]), .C1(n3382), .C2(n2814), .A(n3383), .ZN(n3371) );
  NAND2_X1 U3655 ( .A1(n3370), .A2(n3371), .ZN(p10_muxs_out_2__13_) );
  OAI221_X1 U3656 ( .B1(reg4[9]), .B2(A2[5]), .C1(n2814), .C2(A2[4]), .A(n3384), .ZN(n3372) );
  OAI221_X1 U3657 ( .B1(A2[5]), .B2(reg4[10]), .C1(n3382), .C2(n2810), .A(
        n3383), .ZN(n3373) );
  NAND2_X1 U3658 ( .A1(n3372), .A2(n3373), .ZN(p10_muxs_out_2__14_) );
  OAI221_X1 U3659 ( .B1(reg4[10]), .B2(A2[5]), .C1(n2810), .C2(A2[4]), .A(
        n3384), .ZN(n3374) );
  OAI221_X1 U3660 ( .B1(A2[5]), .B2(reg4[11]), .C1(n3382), .C2(n2861), .A(
        n3383), .ZN(n3375) );
  NAND2_X1 U3661 ( .A1(n3374), .A2(n3375), .ZN(p10_muxs_out_2__15_) );
  OAI221_X1 U3662 ( .B1(reg4[11]), .B2(A2[5]), .C1(n2861), .C2(A2[4]), .A(
        n3384), .ZN(n3376) );
  OAI221_X1 U3663 ( .B1(A2[5]), .B2(reg4[12]), .C1(n3382), .C2(n2858), .A(
        n3383), .ZN(n3377) );
  NAND2_X1 U3664 ( .A1(n3376), .A2(n3377), .ZN(p10_muxs_out_2__16_) );
  AOI22_X1 U3665 ( .A1(A2[5]), .A2(n2859), .B1(reg4[13]), .B2(n3382), .ZN(
        n3378) );
  AOI22_X1 U3666 ( .A1(reg4[12]), .A2(A2[4]), .B1(A2[5]), .B2(n2858), .ZN(
        n3379) );
  AOI22_X1 U3667 ( .A1(n3383), .A2(n3378), .B1(n3379), .B2(n3384), .ZN(
        p10_muxs_out_2__17_) );
  AOI21_X1 U3668 ( .B1(A2[4]), .B2(A2[3]), .A(n2859), .ZN(n3380) );
  OAI21_X1 U3669 ( .B1(A2[4]), .B2(A2[3]), .A(n3382), .ZN(n3381) );
  OAI22_X1 U3670 ( .A1(n3380), .A2(n3382), .B1(n2859), .B2(n3381), .ZN(
        p10_muxs_out_2__18_) );
  NAND2_X1 U3671 ( .A1(reg4[0]), .A2(n3418), .ZN(n3386) );
  XNOR2_X1 U3672 ( .A(n3386), .B(n3416), .ZN(p10_muxs_out_3__6_) );
  OAI221_X1 U3673 ( .B1(reg4[0]), .B2(n3416), .C1(n2839), .C2(A2[6]), .A(n3417), .ZN(n3387) );
  OAI221_X1 U3674 ( .B1(n3416), .B2(reg4[1]), .C1(n3415), .C2(
        p10_minus_A_shifted_14_), .A(n3418), .ZN(n3388) );
  NAND2_X1 U3675 ( .A1(n3387), .A2(n3388), .ZN(p10_muxs_out_3__7_) );
  OAI221_X1 U3676 ( .B1(reg4[1]), .B2(n3416), .C1(p10_minus_A_shifted_14_), 
        .C2(A2[6]), .A(n3417), .ZN(n3389) );
  OAI221_X1 U3677 ( .B1(n3416), .B2(reg4[2]), .C1(n3415), .C2(n2821), .A(n3418), .ZN(n3390) );
  NAND2_X1 U3678 ( .A1(n3389), .A2(n3390), .ZN(p10_muxs_out_3__8_) );
  OAI221_X1 U3679 ( .B1(reg4[2]), .B2(n3416), .C1(n2821), .C2(A2[6]), .A(n3417), .ZN(n3391) );
  OAI221_X1 U3680 ( .B1(n3416), .B2(reg4[3]), .C1(n3415), .C2(
        p10_minus_A_shifted_16_), .A(n3418), .ZN(n3392) );
  NAND2_X1 U3681 ( .A1(n3391), .A2(n3392), .ZN(p10_muxs_out_3__9_) );
  OAI221_X1 U3682 ( .B1(reg4[3]), .B2(n3416), .C1(p10_minus_A_shifted_16_), 
        .C2(A2[6]), .A(n3417), .ZN(n3393) );
  OAI221_X1 U3683 ( .B1(n3416), .B2(reg4[4]), .C1(n3415), .C2(n2818), .A(n3418), .ZN(n3394) );
  NAND2_X1 U3684 ( .A1(n3393), .A2(n3394), .ZN(p10_muxs_out_3__10_) );
  OAI221_X1 U3685 ( .B1(reg4[4]), .B2(n3416), .C1(n2818), .C2(A2[6]), .A(n3417), .ZN(n3395) );
  OAI221_X1 U3686 ( .B1(n3416), .B2(reg4[5]), .C1(n3415), .C2(n2813), .A(n3418), .ZN(n3396) );
  NAND2_X1 U3687 ( .A1(n3395), .A2(n3396), .ZN(p10_muxs_out_3__11_) );
  OAI221_X1 U3688 ( .B1(reg4[5]), .B2(n3416), .C1(n2813), .C2(A2[6]), .A(n3417), .ZN(n3397) );
  OAI221_X1 U3689 ( .B1(n3416), .B2(reg4[6]), .C1(n3415), .C2(n2815), .A(n3418), .ZN(n3398) );
  NAND2_X1 U3690 ( .A1(n3397), .A2(n3398), .ZN(p10_muxs_out_3__12_) );
  OAI221_X1 U3691 ( .B1(reg4[6]), .B2(n3416), .C1(n2815), .C2(A2[6]), .A(n3417), .ZN(n3399) );
  OAI221_X1 U3692 ( .B1(n3416), .B2(reg4[7]), .C1(n3415), .C2(n2830), .A(n3418), .ZN(n3400) );
  NAND2_X1 U3693 ( .A1(n3399), .A2(n3400), .ZN(p10_muxs_out_3__13_) );
  OAI221_X1 U3694 ( .B1(reg4[7]), .B2(n3416), .C1(n2830), .C2(A2[6]), .A(n3417), .ZN(n3401) );
  OAI221_X1 U3695 ( .B1(n3416), .B2(reg4[8]), .C1(n3415), .C2(n2832), .A(n3418), .ZN(n3402) );
  NAND2_X1 U3696 ( .A1(n3401), .A2(n3402), .ZN(p10_muxs_out_3__14_) );
  OAI221_X1 U3697 ( .B1(reg4[8]), .B2(n3416), .C1(n2832), .C2(A2[6]), .A(n3417), .ZN(n3403) );
  OAI221_X1 U3698 ( .B1(n3416), .B2(reg4[9]), .C1(n3415), .C2(n2814), .A(n3418), .ZN(n3404) );
  NAND2_X1 U3699 ( .A1(n3403), .A2(n3404), .ZN(p10_muxs_out_3__15_) );
  OAI221_X1 U3700 ( .B1(reg4[9]), .B2(n3416), .C1(n2814), .C2(A2[6]), .A(n3417), .ZN(n3405) );
  OAI221_X1 U3701 ( .B1(n3416), .B2(reg4[10]), .C1(n3415), .C2(n2810), .A(
        n3418), .ZN(n3406) );
  NAND2_X1 U3702 ( .A1(n3405), .A2(n3406), .ZN(p10_muxs_out_3__16_) );
  OAI221_X1 U3703 ( .B1(reg4[10]), .B2(n3416), .C1(n2810), .C2(A2[6]), .A(
        n3417), .ZN(n3407) );
  OAI221_X1 U3704 ( .B1(n3416), .B2(reg4[11]), .C1(n3415), .C2(n2861), .A(
        n3418), .ZN(n3408) );
  NAND2_X1 U3705 ( .A1(n3407), .A2(n3408), .ZN(p10_muxs_out_3__17_) );
  OAI221_X1 U3706 ( .B1(reg4[11]), .B2(n3416), .C1(n2861), .C2(A2[6]), .A(
        n3417), .ZN(n3409) );
  OAI221_X1 U3707 ( .B1(n3416), .B2(reg4[12]), .C1(n3415), .C2(n2858), .A(
        n3418), .ZN(n3410) );
  NAND2_X1 U3708 ( .A1(n3409), .A2(n3410), .ZN(p10_muxs_out_3__18_) );
  OAI221_X1 U3709 ( .B1(reg4[12]), .B2(n3416), .C1(n2858), .C2(A2[6]), .A(
        n3417), .ZN(n3411) );
  OAI221_X1 U3710 ( .B1(n3416), .B2(reg4[13]), .C1(n3415), .C2(n2859), .A(
        n3418), .ZN(n3412) );
  AOI21_X1 U3711 ( .B1(A2[6]), .B2(A2[5]), .A(n2859), .ZN(n3413) );
  OAI21_X1 U3712 ( .B1(A2[6]), .B2(A2[5]), .A(n3415), .ZN(n3414) );
  OAI22_X1 U3713 ( .A1(n3413), .A2(n3415), .B1(n2859), .B2(n3414), .ZN(
        p10_muxs_out_3__20_) );
  XNOR2_X1 U3714 ( .A(n3419), .B(n1902), .ZN(n1899) );
  XOR2_X1 U3715 ( .A(n1903), .B(n1904), .Z(n3419) );
  XOR2_X1 U3716 ( .A(n1382), .B(n3420), .Z(p11_S[58]) );
  XNOR2_X1 U3717 ( .A(n1384), .B(n1385), .ZN(n3420) );
  XNOR2_X1 U3718 ( .A(p10_muxs_out_2__12_), .B(n1926), .ZN(n1902) );
  AOI222_X1 U3719 ( .A1(n1942), .A2(n1943), .B1(n1942), .B2(n1944), .C1(n1943), 
        .C2(n1944), .ZN(n1721) );
  AOI22_X1 U3720 ( .A1(A1[9]), .A2(n1392), .B1(n1393), .B2(n1394), .ZN(n1391)
         );
  XNOR2_X1 U3721 ( .A(n1641), .B(n1644), .ZN(n1390) );
  AOI222_X1 U3722 ( .A1(n1720), .A2(n1721), .B1(n1720), .B2(n1718), .C1(n1721), 
        .C2(n1718), .ZN(p10_C[59]) );
  XNOR2_X1 U3723 ( .A(n1923), .B(n1945), .ZN(n1720) );
  AOI22_X1 U3724 ( .A1(reg2[13]), .A2(n1406), .B1(n1407), .B2(n2860), .ZN(
        n1405) );
  AOI22_X1 U3725 ( .A1(reg2[12]), .A2(n1406), .B1(n1407), .B2(n2863), .ZN(
        n1423) );
  AOI22_X1 U3726 ( .A1(reg2[11]), .A2(n1406), .B1(n1407), .B2(n2862), .ZN(
        n1428) );
  AOI22_X1 U3727 ( .A1(reg2[10]), .A2(n1406), .B1(n1407), .B2(n2833), .ZN(
        n1449) );
  AOI22_X1 U3728 ( .A1(reg2[7]), .A2(n1406), .B1(n1407), .B2(n2831), .ZN(n1488) );
  AOI22_X1 U3729 ( .A1(reg2[8]), .A2(n1406), .B1(n1407), .B2(n2811), .ZN(n1473) );
  AOI222_X1 U3730 ( .A1(n1597), .A2(p11_muxs_out_3__11_), .B1(n1597), .B2(
        n1598), .C1(p11_muxs_out_3__11_), .C2(n1598), .ZN(n1376) );
  AOI22_X1 U3731 ( .A1(reg2[6]), .A2(n1406), .B1(n1407), .B2(n2835), .ZN(n1507) );
  AOI22_X1 U3732 ( .A1(reg2[4]), .A2(n1406), .B1(n1407), .B2(n2817), .ZN(n1551) );
  AOI22_X1 U3733 ( .A1(reg2[5]), .A2(n1406), .B1(n1407), .B2(n2834), .ZN(n1530) );
  XNOR2_X1 U3734 ( .A(n1597), .B(p11_muxs_out_3__11_), .ZN(n1610) );
  AOI22_X1 U3735 ( .A1(reg2[2]), .A2(n1406), .B1(n1407), .B2(n2820), .ZN(n1593) );
  AOI22_X1 U3736 ( .A1(reg2[3]), .A2(n1406), .B1(n1407), .B2(
        p11_minus_A_shifted_16_), .ZN(n1573) );
  AOI22_X1 U3737 ( .A1(reg2[1]), .A2(n1406), .B1(n1407), .B2(
        p11_minus_A_shifted_14_), .ZN(n1612) );
  NAND2_X1 U3738 ( .A1(n3421), .A2(n1421), .ZN(n1645) );
  XNOR2_X1 U3739 ( .A(p10_muxs_out_2__8_), .B(p10_muxs_out_1__8_), .ZN(n1986)
         );
  AOI222_X1 U3740 ( .A1(p10_muxs_out_2__12_), .A2(p10_muxs_out_3__12_), .B1(
        p10_muxs_out_2__12_), .B2(n1920), .C1(p10_muxs_out_3__12_), .C2(n1920), 
        .ZN(n1878) );
  OAI221_X1 U3741 ( .B1(reg4[3]), .B2(n1760), .C1(p10_minus_A_shifted_16_), 
        .C2(n1761), .A(n1927), .ZN(n1920) );
  NOR2_X1 U3742 ( .A1(n3422), .A2(n1980), .ZN(n1983) );
  XNOR2_X1 U3743 ( .A(n1983), .B(n1988), .ZN(n1736) );
  XNOR2_X1 U3744 ( .A(n1959), .B(n1956), .ZN(n1943) );
  AOI22_X1 U3745 ( .A1(p10_muxs_out_2__10_), .A2(p10_muxs_out_3__10_), .B1(
        n1955), .B2(n1954), .ZN(n1959) );
  XNOR2_X1 U3746 ( .A(p11_muxs_out_2__8_), .B(p11_muxs_out_1__8_), .ZN(n1646)
         );
  XNOR2_X1 U3747 ( .A(n1646), .B(n1631), .ZN(n1641) );
  XOR2_X1 U3748 ( .A(n1560), .B(n3423), .Z(n1377) );
  XNOR2_X1 U3749 ( .A(n1558), .B(n1559), .ZN(n3423) );
  AOI222_X1 U3750 ( .A1(n1602), .A2(n1603), .B1(n1602), .B2(n1604), .C1(n1603), 
        .C2(n1604), .ZN(n1381) );
  NAND2_X1 U3751 ( .A1(p11_muxs_out_3__8_), .A2(n1638), .ZN(n1389) );
  OAI221_X1 U3752 ( .B1(n1632), .B2(n2838), .C1(n1633), .C2(reg2[0]), .A(n1420), .ZN(n1638) );
  NAND2_X1 U3753 ( .A1(p10_muxs_out_3__8_), .A2(n1978), .ZN(n1729) );
  OAI221_X1 U3754 ( .B1(n1972), .B2(n2839), .C1(n1973), .C2(reg4[0]), .A(n1760), .ZN(n1978) );
  AOI22_X1 U3755 ( .A1(reg2[13]), .A2(n1549), .B1(A1[1]), .B2(n2860), .ZN(
        n1533) );
  AOI221_X1 U3756 ( .B1(reg2[9]), .B2(n1549), .C1(n2816), .C2(n1569), .A(n1637), .ZN(n1625) );
  AOI22_X1 U3757 ( .A1(reg2[13]), .A2(n1549), .B1(n1569), .B2(n2860), .ZN(
        n1568) );
  AOI22_X1 U3758 ( .A1(n1608), .A2(n2833), .B1(n1549), .B2(reg2[11]), .ZN(
        n1607) );
  AOI22_X1 U3759 ( .A1(reg2[8]), .A2(n1549), .B1(n1569), .B2(n2811), .ZN(n1647) );
  AOI221_X1 U3760 ( .B1(reg2[6]), .B2(n1549), .C1(n2835), .C2(n1569), .A(n1656), .ZN(n1649) );
  AOI22_X1 U3761 ( .A1(n1608), .A2(n2816), .B1(n1549), .B2(reg2[10]), .ZN(
        n1621) );
  XOR2_X1 U3762 ( .A(n1944), .B(n3425), .Z(n1725) );
  XNOR2_X1 U3763 ( .A(n1942), .B(n1943), .ZN(n3425) );
  NAND2_X1 U3764 ( .A1(n2043), .A2(n3426), .ZN(n2431) );
  XNOR2_X1 U3765 ( .A(n724), .B(n725), .ZN(p7_S[59]) );
  AOI222_X1 U3766 ( .A1(n730), .A2(n731), .B1(n730), .B2(n728), .C1(n731), 
        .C2(n728), .ZN(p7_C[58]) );
  XNOR2_X1 U3767 ( .A(n732), .B(n733), .ZN(p7_S[57]) );
  AOI222_X1 U3768 ( .A1(n736), .A2(n2812), .B1(n736), .B2(n739), .C1(n2812), 
        .C2(n739), .ZN(p7_C[56]) );
  NAND2_X1 U3769 ( .A1(n2012), .A2(n3427), .ZN(n2398) );
  XNOR2_X1 U3770 ( .A(n72), .B(n73), .ZN(p9_S[59]) );
  XNOR2_X1 U3771 ( .A(n80), .B(n81), .ZN(p9_S[57]) );
  AOI222_X1 U3772 ( .A1(n84), .A2(n2789), .B1(n84), .B2(n87), .C1(n2789), .C2(
        n87), .ZN(p9_C[56]) );
  NAND2_X1 U3773 ( .A1(n3428), .A2(n2028), .ZN(n2415) );
  XNOR2_X1 U3774 ( .A(n398), .B(n399), .ZN(p8_S[59]) );
  AOI222_X1 U3775 ( .A1(n404), .A2(n405), .B1(n404), .B2(n402), .C1(n405), 
        .C2(n402), .ZN(p8_C[58]) );
  XNOR2_X1 U3776 ( .A(n406), .B(n407), .ZN(p8_S[57]) );
  AOI222_X1 U3777 ( .A1(n410), .A2(n2788), .B1(n410), .B2(n413), .C1(n2788), 
        .C2(n413), .ZN(p8_C[56]) );
  XNOR2_X1 U3778 ( .A(n978), .B(n983), .ZN(n742) );
  XNOR2_X1 U3779 ( .A(n326), .B(n331), .ZN(n90) );
  XNOR2_X1 U3780 ( .A(n652), .B(n657), .ZN(n416) );
  XNOR2_X1 U3781 ( .A(n1619), .B(n1616), .ZN(n1603) );
  AOI22_X1 U3782 ( .A1(p11_muxs_out_2__10_), .A2(p11_muxs_out_3__10_), .B1(
        n1615), .B2(n1614), .ZN(n1619) );
  XOR2_X1 U3783 ( .A(n1604), .B(n3429), .Z(n1385) );
  XNOR2_X1 U3784 ( .A(n1602), .B(n1603), .ZN(n3429) );
  AOI222_X1 U3785 ( .A1(n1716), .A2(n1717), .B1(n1716), .B2(n1714), .C1(n1717), 
        .C2(n1714), .ZN(p10_C[60]) );
  AOI222_X1 U3786 ( .A1(n1898), .A2(n1899), .B1(n1898), .B2(n1900), .C1(n1899), 
        .C2(n1900), .ZN(n1713) );
  XNOR2_X1 U3787 ( .A(n1730), .B(n1731), .ZN(p10_S[56]) );
  AOI22_X1 U3788 ( .A1(reg4[13]), .A2(n1889), .B1(A2[1]), .B2(n2859), .ZN(
        n1873) );
  AOI221_X1 U3789 ( .B1(reg4[9]), .B2(n1889), .C1(n2814), .C2(n1909), .A(n1977), .ZN(n1965) );
  AOI22_X1 U3790 ( .A1(reg4[13]), .A2(n1889), .B1(n1909), .B2(n2859), .ZN(
        n1908) );
  AOI22_X1 U3791 ( .A1(n1948), .A2(n2810), .B1(n1889), .B2(reg4[11]), .ZN(
        n1947) );
  AOI22_X1 U3792 ( .A1(reg4[8]), .A2(n1889), .B1(n1909), .B2(n2832), .ZN(n1987) );
  AOI221_X1 U3793 ( .B1(reg4[6]), .B2(n1889), .C1(n2815), .C2(n1909), .A(n1996), .ZN(n1989) );
  AOI22_X1 U3794 ( .A1(n1948), .A2(n2814), .B1(n1889), .B2(reg4[10]), .ZN(
        n1961) );
  AOI222_X1 U3795 ( .A1(n1062), .A2(n2819), .B1(n1062), .B2(n1065), .C1(n2819), 
        .C2(n1065), .ZN(p6_C[56]) );
  AOI22_X1 U3796 ( .A1(reg1_reg[9]), .A2(n1064), .B1(n1065), .B2(n2819), .ZN(
        n1063) );
  XOR2_X1 U3797 ( .A(n1722), .B(n3430), .Z(p10_S[58]) );
  XNOR2_X1 U3798 ( .A(n1724), .B(n1725), .ZN(n3430) );
  XNOR2_X1 U3799 ( .A(n1390), .B(n1391), .ZN(p11_S[56]) );
  XNOR2_X1 U3800 ( .A(n1643), .B(n1648), .ZN(n1396) );
  OAI21_X1 U3801 ( .B1(A1[8]), .B2(A1[7]), .A(n1421), .ZN(n3432) );
  OAI21_X1 U3802 ( .B1(A1[8]), .B2(A1[7]), .A(n1421), .ZN(n3431) );
  MUX2_X1 U3803 ( .A(temp6[13]), .B(reg7[13]), .S(n3435), .Z(n2566) );
  XNOR2_X1 U3804 ( .A(n1375), .B(n1374), .ZN(p11_S[60]) );
  AOI222_X1 U3805 ( .A1(n1376), .A2(n1377), .B1(n1376), .B2(n1374), .C1(n1377), 
        .C2(n1374), .ZN(p11_C[60]) );
  OAI21_X1 U3806 ( .B1(A2[8]), .B2(A2[7]), .A(n1761), .ZN(n3434) );
  OAI21_X1 U3807 ( .B1(A2[8]), .B2(A2[7]), .A(n1761), .ZN(n3433) );
  OAI21_X1 U3808 ( .B1(A2[8]), .B2(A2[7]), .A(n1761), .ZN(n1985) );
  NAND2_X1 U3809 ( .A1(VIN), .A2(temp2[13]), .ZN(n2043) );
  AOI21_X1 U3810 ( .B1(n986), .B2(n2855), .A(n975), .ZN(n978) );
  NAND2_X1 U3811 ( .A1(VIN), .A2(temp3[13]), .ZN(n2028) );
  AOI21_X1 U3812 ( .B1(n660), .B2(n2856), .A(n649), .ZN(n652) );
  NAND2_X1 U3813 ( .A1(VIN), .A2(temp4[13]), .ZN(n2012) );
  AOI21_X1 U3814 ( .B1(n334), .B2(n2857), .A(n323), .ZN(n326) );
  OAI221_X1 U3815 ( .B1(reg2[3]), .B2(n1420), .C1(p11_minus_A_shifted_16_), 
        .C2(n1421), .A(n1587), .ZN(n1580) );
  AOI222_X1 U3816 ( .A1(p11_muxs_out_2__12_), .A2(p11_muxs_out_3__12_), .B1(
        p11_muxs_out_2__12_), .B2(n1580), .C1(p11_muxs_out_3__12_), .C2(n1580), 
        .ZN(n1538) );
  XNOR2_X1 U3817 ( .A(n1714), .B(n1715), .ZN(p10_S[60]) );
  XNOR2_X1 U3818 ( .A(n1900), .B(n1924), .ZN(n1717) );
  XNOR2_X1 U3819 ( .A(n1378), .B(n1379), .ZN(p11_S[59]) );
  XNOR2_X1 U3820 ( .A(n1386), .B(n1387), .ZN(p11_S[57]) );
  AOI222_X1 U3821 ( .A1(n1390), .A2(n1394), .B1(n1390), .B2(n1393), .C1(n1394), 
        .C2(n1393), .ZN(p11_C[56]) );
  XNOR2_X1 U3822 ( .A(n1718), .B(n1719), .ZN(p10_S[59]) );
  AOI222_X1 U3823 ( .A1(n1724), .A2(n3424), .B1(n1724), .B2(n1722), .C1(n3424), 
        .C2(n1722), .ZN(p10_C[58]) );
  XNOR2_X1 U3824 ( .A(n1726), .B(n1727), .ZN(p10_S[57]) );
  AOI222_X1 U3825 ( .A1(n1730), .A2(n1734), .B1(n1730), .B2(n1733), .C1(n1734), 
        .C2(n1733), .ZN(p10_C[56]) );
  AOI22_X1 U3826 ( .A1(A2[9]), .A2(n1732), .B1(n1733), .B2(n1734), .ZN(n1731)
         );
  AOI22_X1 U3827 ( .A1(reg4[13]), .A2(n1769), .B1(n1770), .B2(n2859), .ZN(
        n1762) );
  AOI22_X1 U3828 ( .A1(reg4[12]), .A2(n1769), .B1(n1770), .B2(n2858), .ZN(
        n1790) );
  AOI22_X1 U3829 ( .A1(reg4[11]), .A2(n1769), .B1(n1770), .B2(n2861), .ZN(
        n1799) );
  AOI22_X1 U3830 ( .A1(reg4[10]), .A2(n1769), .B1(n1770), .B2(n2810), .ZN(
        n1815) );
  AOI22_X1 U3831 ( .A1(reg4[9]), .A2(n1769), .B1(n1770), .B2(n2814), .ZN(n1825) );
  AOI22_X1 U3832 ( .A1(reg4[8]), .A2(n1769), .B1(n1770), .B2(n2832), .ZN(n1840) );
  AOI22_X1 U3833 ( .A1(reg4[7]), .A2(n1769), .B1(n1770), .B2(n2830), .ZN(n1867) );
  AOI22_X1 U3834 ( .A1(reg4[6]), .A2(n1769), .B1(n1770), .B2(n2815), .ZN(n1888) );
  AOI22_X1 U3835 ( .A1(reg4[3]), .A2(n1769), .B1(n1770), .B2(
        p10_minus_A_shifted_16_), .ZN(n1951) );
  AOI22_X1 U3836 ( .A1(reg4[5]), .A2(n1769), .B1(n1770), .B2(n2813), .ZN(n1911) );
  AOI22_X1 U3837 ( .A1(reg4[2]), .A2(n1769), .B1(n1770), .B2(n2821), .ZN(n1962) );
  AOI22_X1 U3838 ( .A1(reg4[4]), .A2(n1769), .B1(n1770), .B2(n2818), .ZN(n1927) );
  AOI22_X1 U3839 ( .A1(reg2[13]), .A2(n1429), .B1(n1430), .B2(n2860), .ZN(
        n1422) );
  AOI22_X1 U3840 ( .A1(reg2[12]), .A2(n1429), .B1(n1430), .B2(n2863), .ZN(
        n1450) );
  AOI22_X1 U3841 ( .A1(reg2[11]), .A2(n1429), .B1(n1430), .B2(n2862), .ZN(
        n1459) );
  AOI22_X1 U3842 ( .A1(reg2[10]), .A2(n1429), .B1(n1430), .B2(n2833), .ZN(
        n1475) );
  AOI22_X1 U3843 ( .A1(reg2[9]), .A2(n1429), .B1(n1430), .B2(n2816), .ZN(n1485) );
  AOI22_X1 U3844 ( .A1(reg2[8]), .A2(n1429), .B1(n1430), .B2(n2811), .ZN(n1500) );
  AOI22_X1 U3845 ( .A1(reg2[7]), .A2(n1429), .B1(n1430), .B2(n2831), .ZN(n1527) );
  AOI22_X1 U3846 ( .A1(reg2[6]), .A2(n1429), .B1(n1430), .B2(n2835), .ZN(n1548) );
  AOI22_X1 U3847 ( .A1(reg2[3]), .A2(n1429), .B1(n1430), .B2(
        p11_minus_A_shifted_16_), .ZN(n1611) );
  AOI22_X1 U3848 ( .A1(reg2[5]), .A2(n1429), .B1(n1430), .B2(n2834), .ZN(n1571) );
  AOI22_X1 U3849 ( .A1(reg2[2]), .A2(n1429), .B1(n1430), .B2(n2820), .ZN(n1622) );
  AOI22_X1 U3850 ( .A1(reg2[4]), .A2(n1429), .B1(n1430), .B2(n2817), .ZN(n1587) );
  MUX2_X1 U3851 ( .A(n3436), .B(n1917), .S(n2859), .Z(p10_final_product1[26])
         );
  MUX2_X1 U3852 ( .A(n2804), .B(n3437), .S(B3[13]), .Z(p9_final_product1[26])
         );
  MUX2_X1 U3853 ( .A(n2805), .B(n3438), .S(B2[13]), .Z(p8_final_product1[26])
         );
  MUX2_X1 U3854 ( .A(n2866), .B(n3439), .S(B1[13]), .Z(p7_final_product1[26])
         );
  MUX2_X1 U3855 ( .A(n3440), .B(n1577), .S(n2860), .Z(p11_final_product1[26])
         );
endmodule

