
module IIR_ADV ( CLK, RST_n, VIN, DIN, B0, B1, B2, B3, A1, A2, VOUT, DOUT );
  input [13:0] DIN;
  input [13:0] B0;
  input [13:0] B1;
  input [13:0] B2;
  input [13:0] B3;
  input [13:0] A1;
  input [13:0] A2;
  output [13:0] DOUT;
  input CLK, RST_n, VIN;
  output VOUT;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, REGISTER_in_n42, REGISTER_in_n41, REGISTER_in_n40,
         REGISTER_in_n39, REGISTER_in_n38, REGISTER_in_n37, REGISTER_in_n36,
         REGISTER_in_n35, REGISTER_in_n34, REGISTER_in_n33, REGISTER_in_n32,
         REGISTER_in_n31, REGISTER_in_n30, REGISTER_in_n29,
         p6_final_product2_25_, p6_final_product2_26_, p6_final_product1_26,
         SUB1_N1, SUB1_N10, SUB1_N11, SUB1_N12, SUB1_N13, SUB1_N2, SUB1_N3,
         SUB1_N4, SUB1_N5, SUB1_N6, SUB1_N7, SUB1_N8, SUB1_N9, REG61_n62,
         REG61_n61, REG61_n60, REG61_n59, REG61_n58, REG61_n57, REG61_n56,
         REG61_n55, REG61_n54, REG61_n53, REG61_n52, REG61_n51, REG61_n50,
         REG61_n49, REG51_n63, REG51_n62, REG51_n61, REG51_n60, REG51_n59,
         REG51_n58, REG51_n57, REG51_n56, REG51_n55, REG51_n54, REG51_n53,
         REG51_n52, REG51_n51, REG51_n50, REG41_n61, REG41_n60, REG41_n59,
         REG41_n58, REG41_n57, REG41_n56, REG41_n55, REG41_n54, REG41_n53,
         REG41_n52, REG41_n51, REG41_n50, REG41_n49, REG41_n48, REG31_n61,
         REG31_n60, REG31_n59, REG31_n58, REG31_n57, REG31_n56, REG31_n55,
         REG31_n54, REG31_n53, REG31_n52, REG31_n51, REG31_n50, REG31_n49,
         REG31_n48, REG21_n61, REG21_n60, REG21_n59, REG21_n58, REG21_n57,
         REG21_n56, REG21_n55, REG21_n54, REG21_n53, REG21_n52, REG21_n51,
         REG21_n50, REG21_n49, REG21_n48, REG11_n61, REG11_n60, REG11_n59,
         REG11_n58, REG11_n57, REG11_n56, REG11_n55, REG11_n54, REG11_n53,
         REG11_n52, REG11_n51, REG11_n50, REG11_n49, REG11_n48,
         REGISTER_out_n75, REGISTER_out_n74, REGISTER_out_n73,
         REGISTER_out_n72, REGISTER_out_n71, REGISTER_out_n70,
         REGISTER_out_n69, REGISTER_out_n68, REGISTER_out_n67,
         REGISTER_out_n66, REGISTER_out_n65, REGISTER_out_n64,
         REGISTER_out_n63, REGISTER_out_n62, REGISTER_out_n61,
         REGISTER_out_n60, REGISTER_out_n59, REGISTER_out_n58,
         REGISTER_out_n57, REGISTER_out_n56, REGISTER_out_n55,
         REGISTER_out_n54, REGISTER_out_n53, REGISTER_out_n52,
         REGISTER_out_n51, REGISTER_out_n50, REGISTER_out_n49,
         REGISTER_out_n48, REG4_1_n62, REG4_1_n61, REG4_1_n60, REG4_1_n59,
         REG4_1_n58, REG4_1_n57, REG4_1_n56, REG4_1_n55, REG4_1_n54,
         REG4_1_n53, REG4_1_n52, REG4_1_n51, REG4_1_n50, REG4_1_n49,
         REGISTER4_n61, REGISTER4_n60, REGISTER4_n59, REGISTER4_n58,
         REGISTER4_n57, REGISTER4_n56, REGISTER4_n55, REGISTER4_n54,
         REGISTER4_n53, REGISTER4_n52, REGISTER4_n50, REGISTER4_n49,
         REGISTER4_n48, REG3_1_n62, REG3_1_n61, REG3_1_n60, REG3_1_n59,
         REG3_1_n58, REG3_1_n57, REG3_1_n56, REG3_1_n55, REG3_1_n54,
         REG3_1_n53, REG3_1_n52, REG3_1_n51, REG3_1_n50, REG3_1_n49,
         REGISTER3_n61, REGISTER3_n60, REGISTER3_n59, REGISTER3_n58,
         REGISTER3_n57, REGISTER3_n56, REGISTER3_n55, REGISTER3_n54,
         REGISTER3_n53, REGISTER3_n52, REGISTER3_n51, REGISTER3_n50,
         REGISTER3_n49, REGISTER3_n48, REG2_1_n62, REG2_1_n61, REG2_1_n60,
         REG2_1_n59, REG2_1_n58, REG2_1_n57, REG2_1_n56, REG2_1_n55,
         REG2_1_n54, REG2_1_n53, REG2_1_n52, REG2_1_n51, REG2_1_n50,
         REG2_1_n49, REGISTER2_n61, REGISTER2_n60, REGISTER2_n59,
         REGISTER2_n58, REGISTER2_n57, REGISTER2_n56, REGISTER2_n55,
         REGISTER2_n54, REGISTER2_n53, REGISTER2_n52, REGISTER2_n51,
         REGISTER2_n50, REGISTER2_n49, REGISTER2_n48, REG1_1_n62, REG1_1_n61,
         REG1_1_n60, REG1_1_n59, REG1_1_n58, REG1_1_n57, REG1_1_n56,
         REG1_1_n55, REG1_1_n54, REG1_1_n53, REG1_1_n52, REG1_1_n51,
         REG1_1_n50, REG1_1_n49, REGISTER1_n61, REGISTER1_n60, REGISTER1_n59,
         REGISTER1_n58, REGISTER1_n57, REGISTER1_n56, REGISTER1_n55,
         REGISTER1_n54, REGISTER1_n53, REGISTER1_n52, REGISTER1_n51,
         REGISTER1_n50, REGISTER1_n49, REGISTER1_n48, p10_final_product2_25_,
         p10_final_product2_26_, \p10/final_product1[0] ,
         p10_final_product1_26, p11_final_product2_25_, p11_final_product2_26_,
         p11_final_product1_26, p9_final_product2_25_, p9_final_product2_26_,
         p9_final_product1_26, p8_final_product2_25_, p8_final_product2_26_,
         p8_final_product1_26, p7_final_product2_25_, p7_final_product2_26_,
         p7_final_product1_26, sig_ff2_9_, sig_ff2_8_, sig_ff2_7_, sig_ff2_6_,
         sig_ff2_5_, sig_ff2_4_, sig_ff2_3_, sig_ff2_2_, sig_ff2_1_,
         sig_ff2_13_, sig_ff2_12_, sig_ff2_11_, sig_ff2_10_, sig_ff2_0_,
         sig_ff1_9_, sig_ff1_8_, sig_ff1_7_, sig_ff1_6_, sig_ff1_5_,
         sig_ff1_4_, sig_ff1_3_, sig_ff1_2_, sig_ff1_1_, sig_ff1_13_,
         sig_ff1_12_, sig_ff1_11_, sig_ff1_10_, sig_ff1_0_, fb_9_, fb_8_,
         fb_7_, fb_6_, fb_5_, fb_4_, fb_3_, fb_2_, fb_1_, fb_13_, fb_12_,
         fb_11_, fb_10_, fb_0_, n513, n515, n519, n521, n523, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n582, n583, n584,
         n585, n586, n587, n588, n590, n591, n592, n594, n595, n596, n598,
         n599, n600, n602, n603, n604, n605, n606, n607, n608, n609, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n858, n859, n863, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n912, n913, n914, n915, n916, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n972, n973, n975, n976, n977, n978, n979,
         n980, n981, n983, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1040, n1041, n1042, n1044, n1045,
         n1046, n1048, n1049, n1050, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1307, n1308, n1309, n1311, n1313, n1317,
         n1318, n1319, n1320, n1321, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1341, n1342, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1361,
         n1362, n1363, n1364, n1365, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1421, n1422, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1489,
         n1490, n1491, n1493, n1494, n1495, n1497, n1498, n1499, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1757,
         n1758, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1795, n1796, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1811, n1812, n1813, n1814,
         n1815, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1871, n1872, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1940, n1941, n1943, n1944, n1945,
         n1947, n1948, n1949, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1960, n1961, n1962, n1963, n1964, n1965, n1967, n1969, n1970,
         n1971, n1972, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2162, n2163, n2164, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2207, n2208,
         n2212, n2214, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2245, n2246, n2247, n2248,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2261, n2262, n2263, n2264, n2265, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2280, n2281, n2282, n2283, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2304, n2305, n2306, n2307, n2308,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2322, n2324, n2326,
         n2327, n2328, n2329, n2331, n2332, n2333, n2334, n2335, n2337, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2381, n2382, n2383, n2385, n2386, n2387, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2435, n2436, n2437, n2438, n2439, n2440, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2454, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2514, n2515, n2516, n2517, n2518, n2519, n2521,
         n2522, n2523, n2524, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2660, n2661, n2663, n2664, n2666, n2667, n2668, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2685, n2686, n2691, n2692, n2693, n2694, n2695, n2697,
         n2698, n2700, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2766, n2767, n2768, n2769, n2771, n2774,
         n2776, n2777, n2778, n2779, n2781, n2782, n2784, n2785, n2787, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2840, n2841, n2842,
         n2843, n2844, n2845, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2861, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2885, n2886,
         n2887, n2888, n2889, n2890, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2904, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3009, n3010, n3011, n3012, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3105, n3106, n3107, n3109, n3110,
         n3111, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3142, n3143, n3144,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3194, n3195, n3196, n3197,
         n3199, n3200, n3201, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3221,
         n3222, n3224, n3225, n3226, n3228, n3229, n3230, n3231, n3233, n3234,
         n3235, n3236, n3238, n3239, n3240, n3241, n3242, n3244, n3245, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3264, n3266, n3268, n3270, n3272, n3278, n3280,
         n3282, n3284, n3286, n3288, n3290, n3291, n3293, n3294, n3296, n3297,
         n3299, n3300, n3302, n3303, n3305, n3306, n3307, n3308, n3309, n3310,
         n3312, n3313, n3315, n3316, n3318, n3319, n3321, n3322, n3324, n3325,
         n3326, n3327, n1939, n1938, n589, n597, n2846, n1051, n1039, n3202,
         n1496, n1946, n862, n2211, n2659, n1950, n2278, n2266, n1488, n1500,
         n1942, n1312, n1761, n2161,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_,
         SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_, s6_add_23_carry_1_,
         s6_add_23_carry_2_, s6_add_23_carry_3_, s6_add_23_carry_4_,
         s6_add_23_carry_5_, s6_add_23_carry_6_, s6_add_23_carry_7_,
         s6_add_23_carry_8_, s6_add_23_carry_9_, s6_add_23_carry_10_,
         s6_add_23_carry_11_, s6_add_23_carry_12_, s6_add_23_carry_13_,
         s9_add_23_carry_1_, s9_add_23_carry_2_, s9_add_23_carry_3_,
         s9_add_23_carry_4_, s9_add_23_carry_5_, s9_add_23_carry_6_,
         s9_add_23_carry_7_, s9_add_23_carry_8_, s9_add_23_carry_9_,
         s9_add_23_carry_10_, s9_add_23_carry_11_, s9_add_23_carry_12_,
         s9_add_23_carry_13_, s8_add_23_carry_1_, s8_add_23_carry_2_,
         s8_add_23_carry_3_, s8_add_23_carry_4_, s8_add_23_carry_5_,
         s8_add_23_carry_6_, s8_add_23_carry_7_, s8_add_23_carry_8_,
         s8_add_23_carry_9_, s8_add_23_carry_10_, s8_add_23_carry_11_,
         s8_add_23_carry_12_, s8_add_23_carry_13_, s7_add_23_carry_1_,
         s7_add_23_carry_2_, s7_add_23_carry_3_, s7_add_23_carry_4_,
         s7_add_23_carry_5_, s7_add_23_carry_6_, s7_add_23_carry_7_,
         s7_add_23_carry_8_, s7_add_23_carry_9_, s7_add_23_carry_10_,
         s7_add_23_carry_11_, s7_add_23_carry_12_, s7_add_23_carry_13_,
         p6_Partial_products_sum_add_23_n180,
         p6_Partial_products_sum_add_23_n233,
         p6_Partial_products_sum_add_23_n232,
         p6_Partial_products_sum_add_23_n231,
         p6_Partial_products_sum_add_23_n230,
         p6_Partial_products_sum_add_23_n229,
         p6_Partial_products_sum_add_23_n228,
         p6_Partial_products_sum_add_23_n227,
         p6_Partial_products_sum_add_23_n226,
         p6_Partial_products_sum_add_23_n225,
         p6_Partial_products_sum_add_23_n224,
         p6_Partial_products_sum_add_23_n223,
         p6_Partial_products_sum_add_23_n222,
         p6_Partial_products_sum_add_23_n221,
         p6_Partial_products_sum_add_23_n220,
         p6_Partial_products_sum_add_23_n219,
         p6_Partial_products_sum_add_23_n218,
         p6_Partial_products_sum_add_23_n217,
         p6_Partial_products_sum_add_23_n216,
         p6_Partial_products_sum_add_23_n215,
         p6_Partial_products_sum_add_23_n211,
         p6_Partial_products_sum_add_23_n210,
         p6_Partial_products_sum_add_23_n209,
         p6_Partial_products_sum_add_23_n208,
         p6_Partial_products_sum_add_23_n207,
         p6_Partial_products_sum_add_23_n206,
         p6_Partial_products_sum_add_23_n205,
         p6_Partial_products_sum_add_23_n204,
         p6_Partial_products_sum_add_23_n203,
         p6_Partial_products_sum_add_23_n202,
         p6_Partial_products_sum_add_23_n201,
         p6_Partial_products_sum_add_23_n200,
         p6_Partial_products_sum_add_23_n199,
         p6_Partial_products_sum_add_23_n198,
         p6_Partial_products_sum_add_23_n197,
         p6_Partial_products_sum_add_23_n196,
         p6_Partial_products_sum_add_23_n195,
         p6_Partial_products_sum_add_23_n194,
         p6_Partial_products_sum_add_23_n193,
         p6_Partial_products_sum_add_23_n192,
         p6_Partial_products_sum_add_23_n191,
         p6_Partial_products_sum_add_23_n190,
         p6_Partial_products_sum_add_23_n189,
         p6_Partial_products_sum_add_23_n188,
         p6_Partial_products_sum_add_23_n187,
         p6_Partial_products_sum_add_23_n185,
         p6_Partial_products_sum_add_23_n184,
         p6_Partial_products_sum_add_23_n183,
         p6_Partial_products_sum_add_23_n182,
         p6_Partial_products_sum_add_23_n181,
         p6_Partial_products_sum_add_23_n179,
         p6_Partial_products_sum_add_23_n178,
         p6_Partial_products_sum_add_23_n177,
         p6_Partial_products_sum_add_23_n176,
         p6_Partial_products_sum_add_23_n175,
         p6_Partial_products_sum_add_23_n174,
         p10_Partial_products_sum_add_23_n305,
         p10_Partial_products_sum_add_23_n340,
         p10_Partial_products_sum_add_23_n339,
         p10_Partial_products_sum_add_23_n338,
         p10_Partial_products_sum_add_23_n337,
         p10_Partial_products_sum_add_23_n336,
         p10_Partial_products_sum_add_23_n335,
         p10_Partial_products_sum_add_23_n334,
         p10_Partial_products_sum_add_23_n333,
         p10_Partial_products_sum_add_23_n332,
         p10_Partial_products_sum_add_23_n331,
         p10_Partial_products_sum_add_23_n330,
         p10_Partial_products_sum_add_23_n329,
         p10_Partial_products_sum_add_23_n328,
         p10_Partial_products_sum_add_23_n327,
         p10_Partial_products_sum_add_23_n326,
         p10_Partial_products_sum_add_23_n322,
         p10_Partial_products_sum_add_23_n318,
         p10_Partial_products_sum_add_23_n317,
         p10_Partial_products_sum_add_23_n316,
         p10_Partial_products_sum_add_23_n315,
         p10_Partial_products_sum_add_23_n314,
         p10_Partial_products_sum_add_23_n313,
         p10_Partial_products_sum_add_23_n312,
         p10_Partial_products_sum_add_23_n310,
         p10_Partial_products_sum_add_23_n309,
         p10_Partial_products_sum_add_23_n308,
         p10_Partial_products_sum_add_23_n307,
         p10_Partial_products_sum_add_23_n306,
         p10_Partial_products_sum_add_23_n304,
         p10_Partial_products_sum_add_23_n303,
         p10_Partial_products_sum_add_23_n302,
         p10_Partial_products_sum_add_23_n301,
         p10_Partial_products_sum_add_23_n300,
         p10_Partial_products_sum_add_23_n299,
         p10_Partial_products_sum_add_23_n298,
         p10_Partial_products_sum_add_23_n297,
         p10_Partial_products_sum_add_23_n296,
         p10_Partial_products_sum_add_23_n295,
         p10_Partial_products_sum_add_23_n294,
         p10_Partial_products_sum_add_23_n292,
         p10_Partial_products_sum_add_23_n291,
         p10_Partial_products_sum_add_23_n290,
         p10_Partial_products_sum_add_23_n289,
         p10_Partial_products_sum_add_23_n288,
         p10_Partial_products_sum_add_23_n287,
         p10_Partial_products_sum_add_23_n286,
         p10_Partial_products_sum_add_23_n285,
         p10_Partial_products_sum_add_23_n284,
         p10_Partial_products_sum_add_23_n283,
         p10_Partial_products_sum_add_23_n281,
         p10_Partial_products_sum_add_23_n280,
         p10_Partial_products_sum_add_23_n279,
         p10_Partial_products_sum_add_23_n277,
         p11_Partial_products_sum_add_23_n263,
         p11_Partial_products_sum_add_23_n318,
         p11_Partial_products_sum_add_23_n317,
         p11_Partial_products_sum_add_23_n316,
         p11_Partial_products_sum_add_23_n315,
         p11_Partial_products_sum_add_23_n314,
         p11_Partial_products_sum_add_23_n313,
         p11_Partial_products_sum_add_23_n312,
         p11_Partial_products_sum_add_23_n311,
         p11_Partial_products_sum_add_23_n310,
         p11_Partial_products_sum_add_23_n309,
         p11_Partial_products_sum_add_23_n308,
         p11_Partial_products_sum_add_23_n307,
         p11_Partial_products_sum_add_23_n306,
         p11_Partial_products_sum_add_23_n305,
         p11_Partial_products_sum_add_23_n304,
         p11_Partial_products_sum_add_23_n303,
         p11_Partial_products_sum_add_23_n302,
         p11_Partial_products_sum_add_23_n301,
         p11_Partial_products_sum_add_23_n300,
         p11_Partial_products_sum_add_23_n299,
         p11_Partial_products_sum_add_23_n298,
         p11_Partial_products_sum_add_23_n297,
         p11_Partial_products_sum_add_23_n296,
         p11_Partial_products_sum_add_23_n295,
         p11_Partial_products_sum_add_23_n294,
         p11_Partial_products_sum_add_23_n293,
         p11_Partial_products_sum_add_23_n292,
         p11_Partial_products_sum_add_23_n291,
         p11_Partial_products_sum_add_23_n290,
         p11_Partial_products_sum_add_23_n289,
         p11_Partial_products_sum_add_23_n288,
         p11_Partial_products_sum_add_23_n287,
         p11_Partial_products_sum_add_23_n286,
         p11_Partial_products_sum_add_23_n285,
         p11_Partial_products_sum_add_23_n284,
         p11_Partial_products_sum_add_23_n283,
         p11_Partial_products_sum_add_23_n281,
         p11_Partial_products_sum_add_23_n280,
         p11_Partial_products_sum_add_23_n279,
         p11_Partial_products_sum_add_23_n278,
         p11_Partial_products_sum_add_23_n277,
         p11_Partial_products_sum_add_23_n276,
         p11_Partial_products_sum_add_23_n275,
         p11_Partial_products_sum_add_23_n274,
         p11_Partial_products_sum_add_23_n273,
         p11_Partial_products_sum_add_23_n272,
         p11_Partial_products_sum_add_23_n271,
         p11_Partial_products_sum_add_23_n270,
         p11_Partial_products_sum_add_23_n269,
         p11_Partial_products_sum_add_23_n268,
         p11_Partial_products_sum_add_23_n267,
         p11_Partial_products_sum_add_23_n266,
         p11_Partial_products_sum_add_23_n265,
         p11_Partial_products_sum_add_23_n264,
         p11_Partial_products_sum_add_23_n262,
         p11_Partial_products_sum_add_23_n261,
         p11_Partial_products_sum_add_23_n260,
         p11_Partial_products_sum_add_23_n259,
         p11_Partial_products_sum_add_23_n258,
         p9_Partial_products_sum_add_23_n218,
         p9_Partial_products_sum_add_23_n206,
         p9_Partial_products_sum_add_23_n192,
         p9_Partial_products_sum_add_23_n193,
         p9_Partial_products_sum_add_23_n194,
         p9_Partial_products_sum_add_23_n253,
         p9_Partial_products_sum_add_23_n252,
         p9_Partial_products_sum_add_23_n251,
         p9_Partial_products_sum_add_23_n250,
         p9_Partial_products_sum_add_23_n249,
         p9_Partial_products_sum_add_23_n248,
         p9_Partial_products_sum_add_23_n247,
         p9_Partial_products_sum_add_23_n246,
         p9_Partial_products_sum_add_23_n245,
         p9_Partial_products_sum_add_23_n244,
         p9_Partial_products_sum_add_23_n243,
         p9_Partial_products_sum_add_23_n242,
         p9_Partial_products_sum_add_23_n241,
         p9_Partial_products_sum_add_23_n240,
         p9_Partial_products_sum_add_23_n239,
         p9_Partial_products_sum_add_23_n238,
         p9_Partial_products_sum_add_23_n237,
         p9_Partial_products_sum_add_23_n236,
         p9_Partial_products_sum_add_23_n235,
         p9_Partial_products_sum_add_23_n234,
         p9_Partial_products_sum_add_23_n233,
         p9_Partial_products_sum_add_23_n232,
         p9_Partial_products_sum_add_23_n231,
         p9_Partial_products_sum_add_23_n230,
         p9_Partial_products_sum_add_23_n229,
         p9_Partial_products_sum_add_23_n228,
         p9_Partial_products_sum_add_23_n227,
         p9_Partial_products_sum_add_23_n226,
         p9_Partial_products_sum_add_23_n225,
         p9_Partial_products_sum_add_23_n223,
         p9_Partial_products_sum_add_23_n222,
         p9_Partial_products_sum_add_23_n221,
         p9_Partial_products_sum_add_23_n220,
         p9_Partial_products_sum_add_23_n219,
         p9_Partial_products_sum_add_23_n217,
         p9_Partial_products_sum_add_23_n216,
         p9_Partial_products_sum_add_23_n215,
         p9_Partial_products_sum_add_23_n214,
         p9_Partial_products_sum_add_23_n213,
         p9_Partial_products_sum_add_23_n211,
         p9_Partial_products_sum_add_23_n210,
         p9_Partial_products_sum_add_23_n209,
         p9_Partial_products_sum_add_23_n208,
         p9_Partial_products_sum_add_23_n207,
         p9_Partial_products_sum_add_23_n205,
         p9_Partial_products_sum_add_23_n204,
         p9_Partial_products_sum_add_23_n203,
         p9_Partial_products_sum_add_23_n202,
         p9_Partial_products_sum_add_23_n201,
         p9_Partial_products_sum_add_23_n199,
         p9_Partial_products_sum_add_23_n198,
         p9_Partial_products_sum_add_23_n197,
         p9_Partial_products_sum_add_23_n196,
         p8_Partial_products_sum_add_23_n189,
         p8_Partial_products_sum_add_23_n190,
         p8_Partial_products_sum_add_23_n191,
         p8_Partial_products_sum_add_23_n250,
         p8_Partial_products_sum_add_23_n249,
         p8_Partial_products_sum_add_23_n248,
         p8_Partial_products_sum_add_23_n247,
         p8_Partial_products_sum_add_23_n246,
         p8_Partial_products_sum_add_23_n245,
         p8_Partial_products_sum_add_23_n244,
         p8_Partial_products_sum_add_23_n243,
         p8_Partial_products_sum_add_23_n242,
         p8_Partial_products_sum_add_23_n241,
         p8_Partial_products_sum_add_23_n240,
         p8_Partial_products_sum_add_23_n239,
         p8_Partial_products_sum_add_23_n238,
         p8_Partial_products_sum_add_23_n237,
         p8_Partial_products_sum_add_23_n236,
         p8_Partial_products_sum_add_23_n235,
         p8_Partial_products_sum_add_23_n234,
         p8_Partial_products_sum_add_23_n233,
         p8_Partial_products_sum_add_23_n232,
         p8_Partial_products_sum_add_23_n231,
         p8_Partial_products_sum_add_23_n230,
         p8_Partial_products_sum_add_23_n229,
         p8_Partial_products_sum_add_23_n228,
         p8_Partial_products_sum_add_23_n227,
         p8_Partial_products_sum_add_23_n226,
         p8_Partial_products_sum_add_23_n225,
         p8_Partial_products_sum_add_23_n224,
         p8_Partial_products_sum_add_23_n223,
         p8_Partial_products_sum_add_23_n222,
         p8_Partial_products_sum_add_23_n221,
         p8_Partial_products_sum_add_23_n220,
         p8_Partial_products_sum_add_23_n219,
         p8_Partial_products_sum_add_23_n218,
         p8_Partial_products_sum_add_23_n217,
         p8_Partial_products_sum_add_23_n216,
         p8_Partial_products_sum_add_23_n215,
         p8_Partial_products_sum_add_23_n214,
         p8_Partial_products_sum_add_23_n213,
         p8_Partial_products_sum_add_23_n212,
         p8_Partial_products_sum_add_23_n211,
         p8_Partial_products_sum_add_23_n210,
         p8_Partial_products_sum_add_23_n209,
         p8_Partial_products_sum_add_23_n208,
         p8_Partial_products_sum_add_23_n207,
         p8_Partial_products_sum_add_23_n206,
         p8_Partial_products_sum_add_23_n205,
         p8_Partial_products_sum_add_23_n204,
         p8_Partial_products_sum_add_23_n203,
         p8_Partial_products_sum_add_23_n202,
         p8_Partial_products_sum_add_23_n201,
         p8_Partial_products_sum_add_23_n200,
         p8_Partial_products_sum_add_23_n199,
         p8_Partial_products_sum_add_23_n198,
         p8_Partial_products_sum_add_23_n197,
         p8_Partial_products_sum_add_23_n196,
         p8_Partial_products_sum_add_23_n195,
         p8_Partial_products_sum_add_23_n194,
         p8_Partial_products_sum_add_23_n193,
         p7_Partial_products_sum_add_23_n250,
         p7_Partial_products_sum_add_23_n249,
         p7_Partial_products_sum_add_23_n248,
         p7_Partial_products_sum_add_23_n244,
         p7_Partial_products_sum_add_23_n243,
         p7_Partial_products_sum_add_23_n242,
         p7_Partial_products_sum_add_23_n241,
         p7_Partial_products_sum_add_23_n240,
         p7_Partial_products_sum_add_23_n239,
         p7_Partial_products_sum_add_23_n238,
         p7_Partial_products_sum_add_23_n237,
         p7_Partial_products_sum_add_23_n236,
         p7_Partial_products_sum_add_23_n235,
         p7_Partial_products_sum_add_23_n234,
         p7_Partial_products_sum_add_23_n233,
         p7_Partial_products_sum_add_23_n232,
         p7_Partial_products_sum_add_23_n231,
         p7_Partial_products_sum_add_23_n230,
         p7_Partial_products_sum_add_23_n229,
         p7_Partial_products_sum_add_23_n228,
         p7_Partial_products_sum_add_23_n227,
         p7_Partial_products_sum_add_23_n226,
         p7_Partial_products_sum_add_23_n225,
         p7_Partial_products_sum_add_23_n224,
         p7_Partial_products_sum_add_23_n223,
         p7_Partial_products_sum_add_23_n222,
         p7_Partial_products_sum_add_23_n221,
         p7_Partial_products_sum_add_23_n220,
         p7_Partial_products_sum_add_23_n219,
         p7_Partial_products_sum_add_23_n218,
         p7_Partial_products_sum_add_23_n217,
         p7_Partial_products_sum_add_23_n216,
         p7_Partial_products_sum_add_23_n215,
         p7_Partial_products_sum_add_23_n214,
         p7_Partial_products_sum_add_23_n213,
         p7_Partial_products_sum_add_23_n212,
         p7_Partial_products_sum_add_23_n211,
         p7_Partial_products_sum_add_23_n210,
         p7_Partial_products_sum_add_23_n209,
         p7_Partial_products_sum_add_23_n208,
         p7_Partial_products_sum_add_23_n207,
         p7_Partial_products_sum_add_23_n206,
         p7_Partial_products_sum_add_23_n205,
         p7_Partial_products_sum_add_23_n204,
         p7_Partial_products_sum_add_23_n203,
         p7_Partial_products_sum_add_23_n202,
         p7_Partial_products_sum_add_23_n201,
         p7_Partial_products_sum_add_23_n200,
         p7_Partial_products_sum_add_23_n199,
         p7_Partial_products_sum_add_23_n198,
         p7_Partial_products_sum_add_23_n197,
         p7_Partial_products_sum_add_23_n196,
         p7_Partial_products_sum_add_23_n195,
         p7_Partial_products_sum_add_23_n194,
         p7_Partial_products_sum_add_23_n193,
         p7_Partial_products_sum_add_23_n192,
         p7_Partial_products_sum_add_23_n191,
         p7_Partial_products_sum_add_23_n190,
         p7_Partial_products_sum_add_23_n189, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852;
  wire   [13:0] xin_in;
  wire   [13:0] xin;
  wire   [13:0] w;
  wire   [13:0] reg1_reg;
  wire   [13:0] temp1;
  wire   [13:0] mul1_reg;
  wire   [13:0] reg2;
  wire   [13:0] reg2_reg;
  wire   [13:0] temp2;
  wire   [13:0] mul2_reg;
  wire   [13:0] reg3;
  wire   [13:0] reg3_reg;
  wire   [13:0] temp3;
  wire   [13:0] mul3_reg;
  wire   [13:0] reg5;
  wire   [13:0] reg4_reg;
  wire   [13:0] temp4;
  wire   [13:0] mul4_reg;
  wire   [13:0] temp6;
  wire   [13:0] reg4;
  wire   [13:0] temp5;
  wire   [13:0] reg6;
  wire   [13:0] reg7;
  wire   [13:0] ff;
  wire   [54:32] p6_C;
  wire   [54:33] p6_S;
  wire   [54:32] p10_C;
  wire   [54:33] p10_S;
  wire   [0:1] p11_final_product1;
  wire   [54:32] p11_C;
  wire   [54:32] p11_S;
  wire   [54:32] p9_C;
  wire   [54:32] p9_S;
  wire   [54:32] p8_C;
  wire   [54:32] p8_S;
  wire   [0:1] p7_final_product1;
  wire   [54:32] p7_C;
  wire   [54:32] p7_S;

  DFFR_X1 xin_in_reg_13_ ( .D(n45), .CK(CLK), .RN(RST_n), .Q(xin_in[13]) );
  DFFR_X1 xin_in_reg_12_ ( .D(n44), .CK(CLK), .RN(RST_n), .Q(xin_in[12]) );
  DFFR_X1 xin_in_reg_11_ ( .D(n43), .CK(CLK), .RN(RST_n), .Q(xin_in[11]) );
  DFFR_X1 xin_in_reg_10_ ( .D(n42), .CK(CLK), .RN(RST_n), .Q(xin_in[10]) );
  DFFR_X1 xin_in_reg_9_ ( .D(n41), .CK(CLK), .RN(RST_n), .Q(xin_in[9]) );
  DFFR_X1 xin_in_reg_8_ ( .D(n40), .CK(CLK), .RN(RST_n), .Q(xin_in[8]) );
  DFFR_X1 xin_in_reg_7_ ( .D(n39), .CK(CLK), .RN(RST_n), .Q(xin_in[7]) );
  DFFR_X1 xin_in_reg_6_ ( .D(n38), .CK(CLK), .RN(RST_n), .Q(xin_in[6]) );
  DFFR_X1 xin_in_reg_5_ ( .D(n37), .CK(CLK), .RN(RST_n), .Q(xin_in[5]) );
  DFFR_X1 xin_in_reg_4_ ( .D(n36), .CK(CLK), .RN(RST_n), .Q(xin_in[4]) );
  DFFR_X1 xin_in_reg_3_ ( .D(n35), .CK(CLK), .RN(RST_n), .Q(xin_in[3]) );
  DFFR_X1 xin_in_reg_2_ ( .D(n34), .CK(CLK), .RN(RST_n), .Q(xin_in[2]) );
  DFFR_X1 xin_in_reg_1_ ( .D(n33), .CK(CLK), .RN(RST_n), .Q(xin_in[1]) );
  DFFR_X1 xin_in_reg_0_ ( .D(n32), .CK(CLK), .RN(RST_n), .Q(xin_in[0]) );
  DFFR_X1 VOUT_reg ( .D(n31), .CK(CLK), .RN(RST_n), .Q(VOUT), .QN(n30) );
  DFFR_X1 REGISTER_in_q_reg_0_ ( .D(REGISTER_in_n29), .CK(CLK), .RN(RST_n), 
        .Q(xin[0]) );
  DFFR_X1 REGISTER_in_q_reg_1_ ( .D(REGISTER_in_n30), .CK(CLK), .RN(RST_n), 
        .Q(xin[1]) );
  DFFR_X1 REGISTER_in_q_reg_2_ ( .D(REGISTER_in_n31), .CK(CLK), .RN(RST_n), 
        .Q(xin[2]) );
  DFFR_X1 REGISTER_in_q_reg_3_ ( .D(REGISTER_in_n32), .CK(CLK), .RN(RST_n), 
        .Q(xin[3]) );
  DFFR_X1 REGISTER_in_q_reg_4_ ( .D(REGISTER_in_n33), .CK(CLK), .RN(RST_n), 
        .Q(xin[4]) );
  DFFR_X1 REGISTER_in_q_reg_5_ ( .D(REGISTER_in_n34), .CK(CLK), .RN(RST_n), 
        .Q(xin[5]) );
  DFFR_X1 REGISTER_in_q_reg_6_ ( .D(REGISTER_in_n35), .CK(CLK), .RN(RST_n), 
        .Q(xin[6]) );
  DFFR_X1 REGISTER_in_q_reg_7_ ( .D(REGISTER_in_n36), .CK(CLK), .RN(RST_n), 
        .Q(xin[7]) );
  DFFR_X1 REGISTER_in_q_reg_8_ ( .D(REGISTER_in_n37), .CK(CLK), .RN(RST_n), 
        .Q(xin[8]) );
  DFFR_X1 REGISTER_in_q_reg_9_ ( .D(REGISTER_in_n38), .CK(CLK), .RN(RST_n), 
        .Q(xin[9]) );
  DFFR_X1 REGISTER_in_q_reg_10_ ( .D(REGISTER_in_n39), .CK(CLK), .RN(RST_n), 
        .Q(xin[10]) );
  DFFR_X1 REGISTER_in_q_reg_11_ ( .D(REGISTER_in_n40), .CK(CLK), .RN(RST_n), 
        .Q(xin[11]) );
  DFFR_X1 REGISTER_in_q_reg_12_ ( .D(REGISTER_in_n41), .CK(CLK), .RN(RST_n), 
        .Q(xin[12]) );
  DFFR_X1 REGISTER_in_q_reg_13_ ( .D(REGISTER_in_n42), .CK(CLK), .RN(RST_n), 
        .Q(xin[13]) );
  DFFR_X1 REG61_q_reg_0_ ( .D(REG61_n62), .CK(CLK), .RN(RST_n), .Q(reg7[0]), 
        .QN(n3707) );
  DFFR_X1 REG61_q_reg_1_ ( .D(REG61_n61), .CK(CLK), .RN(RST_n), .Q(reg7[1]), 
        .QN(n3731) );
  DFFR_X1 REG61_q_reg_2_ ( .D(REG61_n60), .CK(CLK), .RN(RST_n), .Q(reg7[2]) );
  DFFR_X1 REG61_q_reg_3_ ( .D(REG61_n59), .CK(CLK), .RN(RST_n), .Q(reg7[3]), 
        .QN(n3727) );
  DFFR_X1 REG61_q_reg_4_ ( .D(REG61_n58), .CK(CLK), .RN(RST_n), .Q(reg7[4]) );
  DFFR_X1 REG61_q_reg_5_ ( .D(REG61_n57), .CK(CLK), .RN(RST_n), .Q(reg7[5]), 
        .QN(n3728) );
  DFFR_X1 REG61_q_reg_6_ ( .D(REG61_n56), .CK(CLK), .RN(RST_n), .Q(reg7[6]) );
  DFFR_X1 REG61_q_reg_7_ ( .D(REG61_n55), .CK(CLK), .RN(RST_n), .Q(reg7[7]), 
        .QN(n3729) );
  DFFR_X1 REG61_q_reg_8_ ( .D(REG61_n54), .CK(CLK), .RN(RST_n), .Q(reg7[8]) );
  DFFR_X1 REG61_q_reg_9_ ( .D(REG61_n53), .CK(CLK), .RN(RST_n), .Q(reg7[9]), 
        .QN(n3730) );
  DFFR_X1 REG61_q_reg_10_ ( .D(REG61_n52), .CK(CLK), .RN(RST_n), .Q(reg7[10])
         );
  DFFR_X1 REG61_q_reg_11_ ( .D(REG61_n51), .CK(CLK), .RN(RST_n), .Q(reg7[11]), 
        .QN(n3748) );
  DFFR_X1 REG61_q_reg_12_ ( .D(REG61_n50), .CK(CLK), .RN(RST_n), .Q(reg7[12])
         );
  DFFR_X1 REG61_q_reg_13_ ( .D(REG61_n49), .CK(CLK), .RN(RST_n), .Q(reg7[13])
         );
  DFFR_X1 REG51_q_reg_0_ ( .D(REG51_n63), .CK(CLK), .RN(RST_n), .Q(reg6[0]), 
        .QN(n3466) );
  DFFR_X1 REG51_q_reg_1_ ( .D(REG51_n62), .CK(CLK), .RN(RST_n), .Q(reg6[1]), 
        .QN(n3474) );
  DFFR_X1 REG51_q_reg_2_ ( .D(REG51_n61), .CK(CLK), .RN(RST_n), .Q(reg6[2]), 
        .QN(n3473) );
  DFFR_X1 REG51_q_reg_3_ ( .D(REG51_n60), .CK(CLK), .RN(RST_n), .Q(reg6[3]), 
        .QN(n3472) );
  DFFR_X1 REG51_q_reg_4_ ( .D(REG51_n59), .CK(CLK), .RN(RST_n), .Q(reg6[4]), 
        .QN(n3471) );
  DFFR_X1 REG51_q_reg_5_ ( .D(REG51_n58), .CK(CLK), .RN(RST_n), .Q(reg6[5]), 
        .QN(n3470) );
  DFFR_X1 REG51_q_reg_6_ ( .D(REG51_n57), .CK(CLK), .RN(RST_n), .Q(reg6[6]), 
        .QN(n3469) );
  DFFR_X1 REG51_q_reg_7_ ( .D(REG51_n56), .CK(CLK), .RN(RST_n), .Q(reg6[7]), 
        .QN(n3468) );
  DFFR_X1 REG51_q_reg_8_ ( .D(REG51_n55), .CK(CLK), .RN(RST_n), .Q(reg6[8]), 
        .QN(n3467) );
  DFFR_X1 REG51_q_reg_9_ ( .D(REG51_n54), .CK(CLK), .RN(RST_n), .Q(reg6[9]), 
        .QN(n3479) );
  DFFR_X1 REG51_q_reg_10_ ( .D(REG51_n53), .CK(CLK), .RN(RST_n), .Q(reg6[10]), 
        .QN(n3478) );
  DFFR_X1 REG51_q_reg_11_ ( .D(REG51_n52), .CK(CLK), .RN(RST_n), .Q(reg6[11]), 
        .QN(n3477) );
  DFFR_X1 REG51_q_reg_12_ ( .D(REG51_n51), .CK(CLK), .RN(RST_n), .Q(reg6[12]), 
        .QN(n3476) );
  DFFR_X1 REG51_q_reg_13_ ( .D(REG51_n50), .CK(CLK), .RN(RST_n), .Q(reg6[13]), 
        .QN(n3475) );
  DFFR_X1 REG41_q_reg_0_ ( .D(REG41_n61), .CK(CLK), .RN(RST_n), .QN(n3747) );
  DFFR_X1 REG41_q_reg_1_ ( .D(REG41_n60), .CK(CLK), .RN(RST_n), .QN(n3746) );
  DFFR_X1 REG41_q_reg_2_ ( .D(REG41_n59), .CK(CLK), .RN(RST_n), .Q(reg5[2]), 
        .QN(n3772) );
  DFFR_X1 REG41_q_reg_3_ ( .D(REG41_n58), .CK(CLK), .RN(RST_n), .QN(n3745) );
  DFFR_X1 REG41_q_reg_4_ ( .D(REG41_n57), .CK(CLK), .RN(RST_n), .Q(reg5[4]), 
        .QN(n3771) );
  DFFR_X1 REG41_q_reg_5_ ( .D(REG41_n56), .CK(CLK), .RN(RST_n), .QN(n3744) );
  DFFR_X1 REG41_q_reg_6_ ( .D(REG41_n55), .CK(CLK), .RN(RST_n), .Q(reg5[6]), 
        .QN(n3770) );
  DFFR_X1 REG41_q_reg_7_ ( .D(REG41_n54), .CK(CLK), .RN(RST_n), .QN(n3743) );
  DFFR_X1 REG41_q_reg_8_ ( .D(REG41_n53), .CK(CLK), .RN(RST_n), .Q(reg5[8]), 
        .QN(n3769) );
  DFFR_X1 REG41_q_reg_9_ ( .D(REG41_n52), .CK(CLK), .RN(RST_n), .QN(n3742) );
  DFFR_X1 REG41_q_reg_10_ ( .D(REG41_n51), .CK(CLK), .RN(RST_n), .Q(reg5[10]), 
        .QN(n3768) );
  DFFR_X1 REG41_q_reg_11_ ( .D(REG41_n50), .CK(CLK), .RN(RST_n), .QN(n3741) );
  DFFR_X1 REG41_q_reg_12_ ( .D(REG41_n49), .CK(CLK), .RN(RST_n), .QN(n3740) );
  DFFR_X1 REG41_q_reg_13_ ( .D(REG41_n48), .CK(CLK), .RN(RST_n), .QN(n3739) );
  DFFR_X1 REG31_q_reg_1_ ( .D(REG31_n60), .CK(CLK), .RN(RST_n), .Q(reg4[1]), 
        .QN(n3666) );
  DFFR_X1 REG31_q_reg_2_ ( .D(REG31_n59), .CK(CLK), .RN(RST_n), .Q(reg4[2]), 
        .QN(n3673) );
  DFFR_X1 REG31_q_reg_3_ ( .D(REG31_n58), .CK(CLK), .RN(RST_n), .Q(reg4[3]), 
        .QN(n3665) );
  DFFR_X1 REG31_q_reg_4_ ( .D(REG31_n57), .CK(CLK), .RN(RST_n), .Q(reg4[4]), 
        .QN(n3668) );
  DFFR_X1 REG31_q_reg_5_ ( .D(REG31_n56), .CK(CLK), .RN(RST_n), .Q(reg4[5]), 
        .QN(n3664) );
  DFFR_X1 REG31_q_reg_7_ ( .D(REG31_n54), .CK(CLK), .RN(RST_n), .Q(reg4[7]), 
        .QN(n3672) );
  DFFR_X1 REG31_q_reg_8_ ( .D(REG31_n53), .CK(CLK), .RN(RST_n), .Q(reg4[8]), 
        .QN(n3667) );
  DFFR_X1 REG31_q_reg_10_ ( .D(REG31_n51), .CK(CLK), .RN(RST_n), .Q(reg4[10]), 
        .QN(n3682) );
  DFFR_X1 REG31_q_reg_11_ ( .D(REG31_n50), .CK(CLK), .RN(RST_n), .Q(reg4[11]), 
        .QN(n3671) );
  DFFR_X1 REG31_q_reg_12_ ( .D(REG31_n49), .CK(CLK), .RN(RST_n), .Q(reg4[12]), 
        .QN(n3679) );
  DFFR_X1 REG31_q_reg_13_ ( .D(REG31_n48), .CK(CLK), .RN(RST_n), .Q(reg4[13]), 
        .QN(n3676) );
  DFFR_X1 REG21_q_reg_0_ ( .D(REG21_n61), .CK(CLK), .RN(RST_n), .QN(n3738) );
  DFFR_X1 REG21_q_reg_1_ ( .D(REG21_n60), .CK(CLK), .RN(RST_n), .QN(n3737) );
  DFFR_X1 REG21_q_reg_2_ ( .D(REG21_n59), .CK(CLK), .RN(RST_n), .Q(reg3[2]), 
        .QN(n3767) );
  DFFR_X1 REG21_q_reg_3_ ( .D(REG21_n58), .CK(CLK), .RN(RST_n), .QN(n3736) );
  DFFR_X1 REG21_q_reg_4_ ( .D(REG21_n57), .CK(CLK), .RN(RST_n), .Q(reg3[4]), 
        .QN(n3766) );
  DFFR_X1 REG21_q_reg_5_ ( .D(REG21_n56), .CK(CLK), .RN(RST_n), .QN(n3735) );
  DFFR_X1 REG21_q_reg_6_ ( .D(REG21_n55), .CK(CLK), .RN(RST_n), .Q(reg3[6]), 
        .QN(n3765) );
  DFFR_X1 REG21_q_reg_7_ ( .D(REG21_n54), .CK(CLK), .RN(RST_n), .QN(n3734) );
  DFFR_X1 REG21_q_reg_8_ ( .D(REG21_n53), .CK(CLK), .RN(RST_n), .Q(reg3[8]), 
        .QN(n3764) );
  DFFR_X1 REG21_q_reg_9_ ( .D(REG21_n52), .CK(CLK), .RN(RST_n), .QN(n3733) );
  DFFR_X1 REG21_q_reg_10_ ( .D(REG21_n51), .CK(CLK), .RN(RST_n), .Q(reg3[10]), 
        .QN(n3763) );
  DFFR_X1 REG21_q_reg_11_ ( .D(REG21_n50), .CK(CLK), .RN(RST_n), .QN(n3732) );
  DFFR_X1 REG21_q_reg_12_ ( .D(REG21_n49), .CK(CLK), .RN(RST_n), .Q(reg3[12]), 
        .QN(n3762) );
  DFFR_X1 REG21_q_reg_13_ ( .D(REG21_n48), .CK(CLK), .RN(RST_n), .QN(n3708) );
  DFFR_X1 REG11_q_reg_2_ ( .D(REG11_n59), .CK(CLK), .RN(RST_n), .Q(reg2[2]), 
        .QN(n3692) );
  DFFR_X1 REG11_q_reg_0_ ( .D(REG11_n61), .CK(CLK), .RN(RST_n), .Q(reg2[0]), 
        .QN(n3689) );
  DFFR_X1 REG11_q_reg_1_ ( .D(REG11_n60), .CK(CLK), .RN(RST_n), .Q(reg2[1]), 
        .QN(n3684) );
  DFFR_X1 REG11_q_reg_3_ ( .D(REG11_n58), .CK(CLK), .RN(RST_n), .Q(reg2[3]), 
        .QN(n3669) );
  DFFR_X1 REG11_q_reg_5_ ( .D(REG11_n56), .CK(CLK), .RN(RST_n), .Q(reg2[5]), 
        .QN(n3677) );
  DFFR_X1 REG11_q_reg_10_ ( .D(REG11_n51), .CK(CLK), .RN(RST_n), .Q(reg2[10]), 
        .QN(n3693) );
  DFFR_X1 REG11_q_reg_13_ ( .D(REG11_n48), .CK(CLK), .RN(RST_n), .Q(reg2[13]), 
        .QN(n3680) );
  DFFR_X1 REGISTER_out_q_reg_0_ ( .D(REGISTER_out_n61), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[0]), .QN(REGISTER_out_n62) );
  DFFR_X1 REGISTER_out_q_reg_1_ ( .D(REGISTER_out_n60), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[1]), .QN(REGISTER_out_n63) );
  DFFR_X1 REGISTER_out_q_reg_2_ ( .D(REGISTER_out_n59), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[2]), .QN(REGISTER_out_n64) );
  DFFR_X1 REGISTER_out_q_reg_3_ ( .D(REGISTER_out_n58), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[3]), .QN(REGISTER_out_n65) );
  DFFR_X1 REGISTER_out_q_reg_4_ ( .D(REGISTER_out_n57), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[4]), .QN(REGISTER_out_n66) );
  DFFR_X1 REGISTER_out_q_reg_5_ ( .D(REGISTER_out_n56), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[5]), .QN(REGISTER_out_n67) );
  DFFR_X1 REGISTER_out_q_reg_6_ ( .D(REGISTER_out_n55), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[6]), .QN(REGISTER_out_n68) );
  DFFR_X1 REGISTER_out_q_reg_7_ ( .D(REGISTER_out_n54), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[7]), .QN(REGISTER_out_n69) );
  DFFR_X1 REGISTER_out_q_reg_8_ ( .D(REGISTER_out_n53), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[8]), .QN(REGISTER_out_n70) );
  DFFR_X1 REGISTER_out_q_reg_9_ ( .D(REGISTER_out_n52), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[9]), .QN(REGISTER_out_n71) );
  DFFR_X1 REGISTER_out_q_reg_10_ ( .D(REGISTER_out_n51), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[10]), .QN(REGISTER_out_n72) );
  DFFR_X1 REGISTER_out_q_reg_11_ ( .D(REGISTER_out_n50), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[11]), .QN(REGISTER_out_n73) );
  DFFR_X1 REGISTER_out_q_reg_12_ ( .D(REGISTER_out_n49), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[12]), .QN(REGISTER_out_n74) );
  DFFR_X1 REGISTER_out_q_reg_13_ ( .D(REGISTER_out_n48), .CK(CLK), .RN(RST_n), 
        .Q(DOUT[13]), .QN(REGISTER_out_n75) );
  DFFR_X1 REG4_1_q_reg_0_ ( .D(REG4_1_n62), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[0]) );
  DFFR_X1 REG4_1_q_reg_1_ ( .D(REG4_1_n61), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[1]) );
  DFFR_X1 REG4_1_q_reg_2_ ( .D(REG4_1_n60), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[2]) );
  DFFR_X1 REG4_1_q_reg_3_ ( .D(REG4_1_n59), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[3]) );
  DFFR_X1 REG4_1_q_reg_4_ ( .D(REG4_1_n58), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[4]) );
  DFFR_X1 REG4_1_q_reg_5_ ( .D(REG4_1_n57), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[5]) );
  DFFR_X1 REG4_1_q_reg_6_ ( .D(REG4_1_n56), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[6]) );
  DFFR_X1 REG4_1_q_reg_7_ ( .D(REG4_1_n55), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[7]) );
  DFFR_X1 REG4_1_q_reg_8_ ( .D(REG4_1_n54), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[8]) );
  DFFR_X1 REG4_1_q_reg_9_ ( .D(REG4_1_n53), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[9]) );
  DFFR_X1 REG4_1_q_reg_10_ ( .D(REG4_1_n52), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[10]) );
  DFFR_X1 REG4_1_q_reg_11_ ( .D(REG4_1_n51), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[11]) );
  DFFR_X1 REG4_1_q_reg_12_ ( .D(REG4_1_n50), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[12]) );
  DFFR_X1 REG4_1_q_reg_13_ ( .D(REG4_1_n49), .CK(CLK), .RN(RST_n), .Q(
        mul4_reg[13]) );
  DFFR_X1 REGISTER4_q_reg_0_ ( .D(REGISTER4_n61), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[0]), .QN(n3705) );
  DFFR_X1 REGISTER4_q_reg_2_ ( .D(REGISTER4_n59), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[2]) );
  DFFR_X1 REGISTER4_q_reg_3_ ( .D(REGISTER4_n58), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[3]), .QN(n3703) );
  DFFR_X1 REGISTER4_q_reg_4_ ( .D(REGISTER4_n57), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[4]) );
  DFFR_X1 REGISTER4_q_reg_5_ ( .D(REGISTER4_n56), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[5]), .QN(n3699) );
  DFFR_X1 REGISTER4_q_reg_6_ ( .D(REGISTER4_n55), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[6]) );
  DFFR_X1 REGISTER4_q_reg_7_ ( .D(REGISTER4_n54), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[7]), .QN(n3697) );
  DFFR_X1 REGISTER4_q_reg_8_ ( .D(REGISTER4_n53), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[8]) );
  DFFR_X1 REGISTER4_q_reg_9_ ( .D(REGISTER4_n52), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[9]), .QN(n3720) );
  DFFR_X1 REGISTER4_q_reg_11_ ( .D(REGISTER4_n50), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[11]), .QN(n3675) );
  DFFR_X1 REGISTER4_q_reg_12_ ( .D(REGISTER4_n49), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[12]), .QN(n3706) );
  DFFR_X1 REG3_1_q_reg_0_ ( .D(REG3_1_n62), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[0]) );
  DFFR_X1 REG3_1_q_reg_1_ ( .D(REG3_1_n61), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[1]) );
  DFFR_X1 REG3_1_q_reg_2_ ( .D(REG3_1_n60), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[2]) );
  DFFR_X1 REG3_1_q_reg_3_ ( .D(REG3_1_n59), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[3]) );
  DFFR_X1 REG3_1_q_reg_4_ ( .D(REG3_1_n58), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[4]) );
  DFFR_X1 REG3_1_q_reg_5_ ( .D(REG3_1_n57), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[5]) );
  DFFR_X1 REG3_1_q_reg_6_ ( .D(REG3_1_n56), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[6]) );
  DFFR_X1 REG3_1_q_reg_7_ ( .D(REG3_1_n55), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[7]) );
  DFFR_X1 REG3_1_q_reg_8_ ( .D(REG3_1_n54), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[8]) );
  DFFR_X1 REG3_1_q_reg_9_ ( .D(REG3_1_n53), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[9]) );
  DFFR_X1 REG3_1_q_reg_10_ ( .D(REG3_1_n52), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[10]) );
  DFFR_X1 REG3_1_q_reg_11_ ( .D(REG3_1_n51), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[11]) );
  DFFR_X1 REG3_1_q_reg_12_ ( .D(REG3_1_n50), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[12]) );
  DFFR_X1 REG3_1_q_reg_13_ ( .D(REG3_1_n49), .CK(CLK), .RN(RST_n), .Q(
        mul3_reg[13]) );
  DFFR_X1 REGISTER3_q_reg_0_ ( .D(REGISTER3_n61), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[0]), .QN(n3704) );
  DFFR_X1 REGISTER3_q_reg_2_ ( .D(REGISTER3_n59), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[2]) );
  DFFR_X1 REGISTER3_q_reg_3_ ( .D(REGISTER3_n58), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[3]), .QN(n3702) );
  DFFR_X1 REGISTER3_q_reg_4_ ( .D(REGISTER3_n57), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[4]) );
  DFFR_X1 REGISTER3_q_reg_5_ ( .D(REGISTER3_n56), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[5]), .QN(n3698) );
  DFFR_X1 REGISTER3_q_reg_6_ ( .D(REGISTER3_n55), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[6]) );
  DFFR_X1 REGISTER3_q_reg_7_ ( .D(REGISTER3_n54), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[7]), .QN(n3696) );
  DFFR_X1 REGISTER3_q_reg_8_ ( .D(REGISTER3_n53), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[8]) );
  DFFR_X1 REGISTER3_q_reg_9_ ( .D(REGISTER3_n52), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[9]), .QN(n3721) );
  DFFR_X1 REGISTER3_q_reg_10_ ( .D(REGISTER3_n51), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[10]) );
  DFFR_X1 REGISTER3_q_reg_11_ ( .D(REGISTER3_n50), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[11]), .QN(n3695) );
  DFFR_X1 REGISTER3_q_reg_12_ ( .D(REGISTER3_n49), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[12]) );
  DFFR_X1 REGISTER3_q_reg_13_ ( .D(REGISTER3_n48), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[13]), .QN(n3761) );
  DFFR_X1 REG2_1_q_reg_0_ ( .D(REG2_1_n62), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[0]) );
  DFFR_X1 REG2_1_q_reg_1_ ( .D(REG2_1_n61), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[1]) );
  DFFR_X1 REG2_1_q_reg_2_ ( .D(REG2_1_n60), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[2]) );
  DFFR_X1 REG2_1_q_reg_3_ ( .D(REG2_1_n59), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[3]) );
  DFFR_X1 REG2_1_q_reg_4_ ( .D(REG2_1_n58), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[4]) );
  DFFR_X1 REG2_1_q_reg_5_ ( .D(REG2_1_n57), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[5]) );
  DFFR_X1 REG2_1_q_reg_6_ ( .D(REG2_1_n56), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[6]) );
  DFFR_X1 REG2_1_q_reg_7_ ( .D(REG2_1_n55), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[7]) );
  DFFR_X1 REG2_1_q_reg_8_ ( .D(REG2_1_n54), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[8]) );
  DFFR_X1 REG2_1_q_reg_9_ ( .D(REG2_1_n53), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[9]) );
  DFFR_X1 REG2_1_q_reg_10_ ( .D(REG2_1_n52), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[10]) );
  DFFR_X1 REG2_1_q_reg_11_ ( .D(REG2_1_n51), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[11]) );
  DFFR_X1 REG2_1_q_reg_12_ ( .D(REG2_1_n50), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[12]) );
  DFFR_X1 REG2_1_q_reg_13_ ( .D(REG2_1_n49), .CK(CLK), .RN(RST_n), .Q(
        mul2_reg[13]) );
  DFFR_X1 REGISTER2_q_reg_0_ ( .D(REGISTER2_n61), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[0]), .QN(n3723) );
  DFFR_X1 REGISTER2_q_reg_2_ ( .D(REGISTER2_n59), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[2]), .QN(n3756) );
  DFFR_X1 REGISTER2_q_reg_4_ ( .D(REGISTER2_n57), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[4]), .QN(n3755) );
  DFFR_X1 REGISTER2_q_reg_5_ ( .D(REGISTER2_n56), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[5]), .QN(n3712) );
  DFFR_X1 REGISTER2_q_reg_6_ ( .D(REGISTER2_n55), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[6]), .QN(n3760) );
  DFFR_X1 REGISTER2_q_reg_7_ ( .D(REGISTER2_n54), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[7]), .QN(n3714) );
  DFFR_X1 REGISTER2_q_reg_8_ ( .D(REGISTER2_n53), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[8]), .QN(n3754) );
  DFFR_X1 REGISTER2_q_reg_9_ ( .D(REGISTER2_n52), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[9]), .QN(n3719) );
  DFFR_X1 REGISTER2_q_reg_10_ ( .D(REGISTER2_n51), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[10]), .QN(n3753) );
  DFFR_X1 REGISTER2_q_reg_11_ ( .D(REGISTER2_n50), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[11]), .QN(n3694) );
  DFFR_X1 REGISTER2_q_reg_12_ ( .D(REGISTER2_n49), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[12]), .QN(n3725) );
  DFFR_X1 REGISTER2_q_reg_13_ ( .D(REGISTER2_n48), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[13]), .QN(n3758) );
  DFFR_X1 REG1_1_q_reg_0_ ( .D(REG1_1_n62), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[0]) );
  DFFR_X1 REG1_1_q_reg_1_ ( .D(REG1_1_n61), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[1]) );
  DFFR_X1 REG1_1_q_reg_2_ ( .D(REG1_1_n60), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[2]) );
  DFFR_X1 REG1_1_q_reg_3_ ( .D(REG1_1_n59), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[3]) );
  DFFR_X1 REG1_1_q_reg_4_ ( .D(REG1_1_n58), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[4]) );
  DFFR_X1 REG1_1_q_reg_5_ ( .D(REG1_1_n57), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[5]) );
  DFFR_X1 REG1_1_q_reg_6_ ( .D(REG1_1_n56), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[6]) );
  DFFR_X1 REG1_1_q_reg_7_ ( .D(REG1_1_n55), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[7]) );
  DFFR_X1 REG1_1_q_reg_8_ ( .D(REG1_1_n54), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[8]) );
  DFFR_X1 REG1_1_q_reg_9_ ( .D(REG1_1_n53), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[9]) );
  DFFR_X1 REG1_1_q_reg_10_ ( .D(REG1_1_n52), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[10]) );
  DFFR_X1 REG1_1_q_reg_11_ ( .D(REG1_1_n51), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[11]) );
  DFFR_X1 REG1_1_q_reg_12_ ( .D(REG1_1_n50), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[12]) );
  DFFR_X1 REG1_1_q_reg_13_ ( .D(REG1_1_n49), .CK(CLK), .RN(RST_n), .Q(
        mul1_reg[13]) );
  DFFR_X1 REGISTER1_q_reg_0_ ( .D(REGISTER1_n61), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[0]), .QN(n3722) );
  DFFR_X1 REGISTER1_q_reg_2_ ( .D(REGISTER1_n59), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[2]), .QN(n3752) );
  DFFR_X1 REGISTER1_q_reg_3_ ( .D(REGISTER1_n58), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[3]), .QN(n3717) );
  DFFR_X1 REGISTER1_q_reg_4_ ( .D(REGISTER1_n57), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[4]), .QN(n3751) );
  DFFR_X1 REGISTER1_q_reg_5_ ( .D(REGISTER1_n56), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[5]), .QN(n3711) );
  DFFR_X1 REGISTER1_q_reg_6_ ( .D(REGISTER1_n55), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[6]), .QN(n3759) );
  DFFR_X1 REGISTER1_q_reg_7_ ( .D(REGISTER1_n54), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[7]), .QN(n3710) );
  DFFR_X1 REGISTER1_q_reg_8_ ( .D(REGISTER1_n53), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[8]), .QN(n3750) );
  DFFR_X1 REGISTER1_q_reg_9_ ( .D(REGISTER1_n52), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[9]), .QN(n3713) );
  DFFR_X1 REGISTER1_q_reg_10_ ( .D(REGISTER1_n51), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[10]), .QN(n3749) );
  DFFR_X1 REGISTER1_q_reg_11_ ( .D(REGISTER1_n50), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[11]), .QN(n3674) );
  DFFR_X1 REGISTER1_q_reg_12_ ( .D(REGISTER1_n49), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[12]), .QN(n3724) );
  DFFR_X1 REGISTER1_q_reg_13_ ( .D(REGISTER1_n48), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[13]), .QN(n3757) );
  MUX2_X1 U2759 ( .A(n3757), .B(n513), .S(B0[13]), .Z(p6_final_product1_26) );
  MUX2_X1 U2760 ( .A(n3758), .B(n515), .S(B1[13]), .Z(p7_final_product1_26) );
  MUX2_X1 U2762 ( .A(n3773), .B(n519), .S(B3[13]), .Z(p9_final_product1_26) );
  MUX2_X1 U2763 ( .A(n521), .B(n2894), .S(n3676), .Z(p10_final_product1_26) );
  MUX2_X1 U2764 ( .A(n523), .B(n2444), .S(n3680), .Z(p11_final_product1_26) );
  XOR2_X1 U2765 ( .A(n543), .B(n544), .Z(n541) );
  XOR2_X1 U2766 ( .A(n550), .B(n551), .Z(n548) );
  XOR2_X1 U2767 ( .A(n554), .B(n555), .Z(n553) );
  XOR2_X1 U2768 ( .A(n558), .B(n559), .Z(n557) );
  XOR2_X1 U2769 ( .A(n562), .B(n563), .Z(n561) );
  XOR2_X1 U2770 ( .A(n566), .B(n567), .Z(n565) );
  XOR2_X1 U2771 ( .A(n570), .B(n571), .Z(n569) );
  XOR2_X1 U2772 ( .A(n574), .B(n575), .Z(n573) );
  XOR2_X1 U2773 ( .A(n576), .B(n577), .Z(p9_S[45]) );
  XOR2_X1 U2775 ( .A(n586), .B(n587), .Z(n585) );
  XOR2_X1 U2781 ( .A(n608), .B(n609), .Z(n607) );
  XOR2_X1 U2782 ( .A(n3697), .B(n611), .Z(p9_S[36]) );
  XOR2_X1 U2783 ( .A(n612), .B(n613), .Z(n611) );
  XOR2_X1 U2784 ( .A(n616), .B(n617), .Z(p9_S[35]) );
  XOR2_X1 U2785 ( .A(n3699), .B(n625), .Z(n622) );
  XOR2_X1 U2786 ( .A(n626), .B(n627), .Z(p9_S[33]) );
  XOR2_X1 U2787 ( .A(n628), .B(n629), .Z(p9_S[32]) );
  XOR2_X1 U2788 ( .A(n3773), .B(n638), .Z(n549) );
  XOR2_X1 U2789 ( .A(n637), .B(n636), .Z(n638) );
  XOR2_X1 U2790 ( .A(n653), .B(n643), .Z(n651) );
  MUX2_X1 U2791 ( .A(n664), .B(n665), .S(n666), .Z(n554) );
  XOR2_X1 U2792 ( .A(n662), .B(n660), .Z(n556) );
  XOR2_X1 U2793 ( .A(n667), .B(n661), .Z(n660) );
  MUX2_X1 U2794 ( .A(n689), .B(n690), .S(n691), .Z(n563) );
  XOR2_X1 U2795 ( .A(n679), .B(n677), .Z(n562) );
  XOR2_X1 U2796 ( .A(n694), .B(n678), .Z(n676) );
  XOR2_X1 U2797 ( .A(n683), .B(n684), .Z(n694) );
  XOR2_X1 U2798 ( .A(n682), .B(n662), .Z(n683) );
  MUX2_X1 U2799 ( .A(n704), .B(n705), .S(n706), .Z(n564) );
  XOR2_X1 U2800 ( .A(n688), .B(n686), .Z(n566) );
  XOR2_X1 U2801 ( .A(n711), .B(n687), .Z(n685) );
  XOR2_X1 U2802 ( .A(n708), .B(n710), .Z(n727) );
  XOR2_X1 U2803 ( .A(n729), .B(n709), .Z(n710) );
  XOR2_X1 U2804 ( .A(n723), .B(n724), .Z(n709) );
  XOR2_X1 U2805 ( .A(n746), .B(n744), .Z(n572) );
  XOR2_X1 U2806 ( .A(n753), .B(n751), .Z(n747) );
  XOR2_X1 U2807 ( .A(n750), .B(n754), .Z(n751) );
  MUX2_X1 U2808 ( .A(n755), .B(n746), .S(n756), .Z(n754) );
  XOR2_X1 U2809 ( .A(n742), .B(n743), .Z(n750) );
  XOR2_X1 U2810 ( .A(n758), .B(n736), .Z(n742) );
  XOR2_X1 U2811 ( .A(n740), .B(n735), .Z(n758) );
  XOR2_X1 U2812 ( .A(n738), .B(n760), .Z(n735) );
  XOR2_X1 U2813 ( .A(n752), .B(n745), .Z(n753) );
  MUX2_X1 U2814 ( .A(n768), .B(n769), .S(n770), .Z(n752) );
  MUX2_X1 U2815 ( .A(n776), .B(n777), .S(n778), .Z(n574) );
  XOR2_X1 U2816 ( .A(n771), .B(n772), .Z(n579) );
  XOR2_X1 U2817 ( .A(n793), .B(n776), .Z(n778) );
  MUX2_X1 U2818 ( .A(n806), .B(n807), .S(n808), .Z(n580) );
  MUX2_X1 U2819 ( .A(n809), .B(n810), .S(n811), .Z(n583) );
  MUX2_X1 U2820 ( .A(n813), .B(n814), .S(n815), .Z(n783) );
  XOR2_X1 U2821 ( .A(n780), .B(n782), .Z(n812) );
  XOR2_X1 U2822 ( .A(n816), .B(n781), .Z(n782) );
  XOR2_X1 U2823 ( .A(n790), .B(n789), .Z(n781) );
  XOR2_X1 U2824 ( .A(n818), .B(n805), .Z(n790) );
  XOR2_X1 U2825 ( .A(n791), .B(n804), .Z(n818) );
  XOR2_X1 U2826 ( .A(n802), .B(n820), .Z(n804) );
  MUX2_X1 U2827 ( .A(n825), .B(n826), .S(n827), .Z(n780) );
  XOR2_X1 U2828 ( .A(n829), .B(n811), .Z(n808) );
  XOR2_X1 U2829 ( .A(n809), .B(n830), .Z(n811) );
  MUX2_X1 U2830 ( .A(n831), .B(n832), .S(n833), .Z(n830) );
  XOR2_X1 U2831 ( .A(n813), .B(n835), .Z(n815) );
  XOR2_X1 U2832 ( .A(n827), .B(n826), .Z(n835) );
  MUX2_X1 U2833 ( .A(n842), .B(n843), .S(n844), .Z(n810) );
  MUX2_X1 U2834 ( .A(n845), .B(n3773), .S(n846), .Z(n587) );
  MUX2_X1 U2835 ( .A(n847), .B(n848), .S(n849), .Z(n586) );
  MUX2_X1 U2836 ( .A(n850), .B(n851), .S(n852), .Z(n588) );
  MUX2_X1 U2837 ( .A(n853), .B(n854), .S(n855), .Z(n591) );
  MUX2_X1 U2841 ( .A(n3675), .B(n874), .S(n875), .Z(n592) );
  MUX2_X1 U2842 ( .A(n876), .B(n877), .S(n878), .Z(n595) );
  XOR2_X1 U2843 ( .A(n852), .B(n851), .Z(n594) );
  XOR2_X1 U2845 ( .A(n898), .B(n876), .Z(n878) );
  XOR2_X1 U2846 ( .A(n884), .B(n885), .Z(n876) );
  MUX2_X1 U2847 ( .A(n904), .B(n905), .S(n906), .Z(n599) );
  MUX2_X1 U2848 ( .A(n907), .B(n908), .S(n909), .Z(n598) );
  MUX2_X1 U2849 ( .A(n910), .B(n3720), .S(n912), .Z(n600) );
  MUX2_X1 U2850 ( .A(n913), .B(n914), .S(n915), .Z(n603) );
  XOR2_X1 U2854 ( .A(n918), .B(n907), .Z(n909) );
  XOR2_X1 U2855 ( .A(n915), .B(n930), .Z(n912) );
  XOR2_X1 U2856 ( .A(n944), .B(n938), .Z(n613) );
  XOR2_X1 U2857 ( .A(n615), .B(n614), .Z(n618) );
  XOR2_X1 U2858 ( .A(n993), .B(n994), .Z(n991) );
  XOR2_X1 U2859 ( .A(n1000), .B(n1001), .Z(n998) );
  XOR2_X1 U2860 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR2_X1 U2861 ( .A(n1008), .B(n1009), .Z(n1007) );
  XOR2_X1 U2862 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR2_X1 U2863 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR2_X1 U2864 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR2_X1 U2865 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR2_X1 U2866 ( .A(n1026), .B(n1027), .Z(p8_S[45]) );
  XOR2_X1 U2867 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR2_X1 U2868 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR2_X1 U2874 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR2_X1 U2875 ( .A(n3696), .B(n1061), .Z(p8_S[36]) );
  XOR2_X1 U2876 ( .A(n1062), .B(n1063), .Z(n1061) );
  XOR2_X1 U2877 ( .A(n1066), .B(n1067), .Z(p8_S[35]) );
  XOR2_X1 U2878 ( .A(n3698), .B(n1075), .Z(n1072) );
  XOR2_X1 U2879 ( .A(n1076), .B(n1077), .Z(p8_S[33]) );
  XOR2_X1 U2880 ( .A(n1078), .B(n1079), .Z(p8_S[32]) );
  XOR2_X1 U2881 ( .A(n3761), .B(n1088), .Z(n999) );
  XOR2_X1 U2882 ( .A(n1087), .B(n1086), .Z(n1088) );
  XOR2_X1 U2883 ( .A(n1103), .B(n1093), .Z(n1101) );
  MUX2_X1 U2884 ( .A(n1114), .B(n1115), .S(n1116), .Z(n1004) );
  XOR2_X1 U2885 ( .A(n1112), .B(n1110), .Z(n1006) );
  XOR2_X1 U2886 ( .A(n1117), .B(n1111), .Z(n1110) );
  MUX2_X1 U2887 ( .A(n1139), .B(n1140), .S(n1141), .Z(n1013) );
  XOR2_X1 U2888 ( .A(n1129), .B(n1127), .Z(n1012) );
  XOR2_X1 U2889 ( .A(n1144), .B(n1128), .Z(n1126) );
  XOR2_X1 U2890 ( .A(n1133), .B(n1134), .Z(n1144) );
  XOR2_X1 U2891 ( .A(n1132), .B(n1112), .Z(n1133) );
  MUX2_X1 U2892 ( .A(n1154), .B(n1155), .S(n1156), .Z(n1014) );
  XOR2_X1 U2893 ( .A(n1138), .B(n1136), .Z(n1016) );
  XOR2_X1 U2894 ( .A(n1161), .B(n1137), .Z(n1135) );
  XOR2_X1 U2895 ( .A(n1158), .B(n1160), .Z(n1177) );
  XOR2_X1 U2896 ( .A(n1179), .B(n1159), .Z(n1160) );
  XOR2_X1 U2897 ( .A(n1173), .B(n1174), .Z(n1159) );
  XOR2_X1 U2898 ( .A(n1196), .B(n1194), .Z(n1022) );
  XOR2_X1 U2899 ( .A(n1203), .B(n1201), .Z(n1197) );
  XOR2_X1 U2900 ( .A(n1200), .B(n1204), .Z(n1201) );
  MUX2_X1 U2901 ( .A(n1205), .B(n1196), .S(n1206), .Z(n1204) );
  XOR2_X1 U2902 ( .A(n1192), .B(n1193), .Z(n1200) );
  XOR2_X1 U2903 ( .A(n1208), .B(n1186), .Z(n1192) );
  XOR2_X1 U2904 ( .A(n1190), .B(n1185), .Z(n1208) );
  XOR2_X1 U2905 ( .A(n1188), .B(n1210), .Z(n1185) );
  XOR2_X1 U2906 ( .A(n1202), .B(n1195), .Z(n1203) );
  MUX2_X1 U2907 ( .A(n1218), .B(n1219), .S(n1220), .Z(n1202) );
  MUX2_X1 U2908 ( .A(n1226), .B(n1227), .S(n1228), .Z(n1024) );
  XOR2_X1 U2909 ( .A(n1221), .B(n1222), .Z(n1029) );
  XOR2_X1 U2910 ( .A(n1243), .B(n1226), .Z(n1228) );
  MUX2_X1 U2911 ( .A(n1256), .B(n1257), .S(n1258), .Z(n1030) );
  MUX2_X1 U2912 ( .A(n1259), .B(n1260), .S(n1261), .Z(n1033) );
  MUX2_X1 U2913 ( .A(n1263), .B(n1264), .S(n1265), .Z(n1233) );
  XOR2_X1 U2914 ( .A(n1230), .B(n1232), .Z(n1262) );
  XOR2_X1 U2915 ( .A(n1266), .B(n1231), .Z(n1232) );
  XOR2_X1 U2916 ( .A(n1240), .B(n1239), .Z(n1231) );
  XOR2_X1 U2917 ( .A(n1268), .B(n1255), .Z(n1240) );
  XOR2_X1 U2918 ( .A(n1241), .B(n1254), .Z(n1268) );
  XOR2_X1 U2919 ( .A(n1252), .B(n1270), .Z(n1254) );
  MUX2_X1 U2920 ( .A(n1275), .B(n1276), .S(n1277), .Z(n1230) );
  XOR2_X1 U2921 ( .A(n1279), .B(n1261), .Z(n1258) );
  XOR2_X1 U2922 ( .A(n1259), .B(n1280), .Z(n1261) );
  MUX2_X1 U2923 ( .A(n1281), .B(n1282), .S(n1283), .Z(n1280) );
  XOR2_X1 U2924 ( .A(n1263), .B(n1285), .Z(n1265) );
  XOR2_X1 U2925 ( .A(n1277), .B(n1276), .Z(n1285) );
  MUX2_X1 U2926 ( .A(n1292), .B(n1293), .S(n1294), .Z(n1260) );
  MUX2_X1 U2927 ( .A(n1295), .B(n3761), .S(n1296), .Z(n1037) );
  MUX2_X1 U2928 ( .A(n1297), .B(n1298), .S(n1299), .Z(n1036) );
  MUX2_X1 U2929 ( .A(n1300), .B(n1301), .S(n1302), .Z(n1038) );
  MUX2_X1 U2930 ( .A(n1303), .B(n1304), .S(n1305), .Z(n1041) );
  MUX2_X1 U2934 ( .A(n3695), .B(n1323), .S(n1324), .Z(n1042) );
  MUX2_X1 U2935 ( .A(n1325), .B(n1326), .S(n1327), .Z(n1045) );
  XOR2_X1 U2937 ( .A(n1344), .B(n1323), .Z(n1324) );
  XOR2_X1 U2938 ( .A(n1347), .B(n1325), .Z(n1327) );
  XOR2_X1 U2939 ( .A(n1333), .B(n1334), .Z(n1325) );
  MUX2_X1 U2940 ( .A(n1353), .B(n1354), .S(n1355), .Z(n1049) );
  MUX2_X1 U2941 ( .A(n1356), .B(n1357), .S(n1358), .Z(n1048) );
  MUX2_X1 U2942 ( .A(n1359), .B(n3721), .S(n1361), .Z(n1050) );
  MUX2_X1 U2943 ( .A(n1362), .B(n1363), .S(n1364), .Z(n1053) );
  XOR2_X1 U2947 ( .A(n1367), .B(n1356), .Z(n1358) );
  XOR2_X1 U2948 ( .A(n1364), .B(n1379), .Z(n1361) );
  XOR2_X1 U2949 ( .A(n1393), .B(n1387), .Z(n1063) );
  XOR2_X1 U2950 ( .A(n1065), .B(n1064), .Z(n1068) );
  XOR2_X1 U2951 ( .A(n1442), .B(n1443), .Z(n1440) );
  XOR2_X1 U2952 ( .A(n1449), .B(n1450), .Z(n1447) );
  XOR2_X1 U2953 ( .A(n1453), .B(n1454), .Z(n1452) );
  XOR2_X1 U2954 ( .A(n1457), .B(n1458), .Z(n1456) );
  XOR2_X1 U2955 ( .A(n1461), .B(n1462), .Z(n1460) );
  XOR2_X1 U2956 ( .A(n1465), .B(n1466), .Z(n1464) );
  XOR2_X1 U2957 ( .A(n1469), .B(n1470), .Z(n1468) );
  XOR2_X1 U2958 ( .A(n1473), .B(n1474), .Z(n1472) );
  XOR2_X1 U2959 ( .A(n1475), .B(n1476), .Z(p7_S[45]) );
  XOR2_X1 U2961 ( .A(n1485), .B(n1486), .Z(n1484) );
  XOR2_X1 U2967 ( .A(n1507), .B(n1508), .Z(n1506) );
  XOR2_X1 U2968 ( .A(n3714), .B(n1510), .Z(p7_S[36]) );
  XOR2_X1 U2969 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR2_X1 U2970 ( .A(n1515), .B(n1516), .Z(p7_S[35]) );
  XOR2_X1 U2971 ( .A(n3712), .B(n1524), .Z(n1521) );
  XOR2_X1 U2972 ( .A(n1525), .B(n1526), .Z(p7_S[33]) );
  XOR2_X1 U2974 ( .A(n3758), .B(n1537), .Z(n1448) );
  XOR2_X1 U2975 ( .A(n1536), .B(n1535), .Z(n1537) );
  XOR2_X1 U2976 ( .A(n1552), .B(n1542), .Z(n1550) );
  MUX2_X1 U2977 ( .A(n1563), .B(n1564), .S(n1565), .Z(n1453) );
  XOR2_X1 U2978 ( .A(n1561), .B(n1559), .Z(n1455) );
  XOR2_X1 U2979 ( .A(n1566), .B(n1560), .Z(n1559) );
  MUX2_X1 U2980 ( .A(n1588), .B(n1589), .S(n1590), .Z(n1462) );
  XOR2_X1 U2981 ( .A(n1578), .B(n1576), .Z(n1461) );
  XOR2_X1 U2982 ( .A(n1593), .B(n1577), .Z(n1575) );
  XOR2_X1 U2983 ( .A(n1582), .B(n1583), .Z(n1593) );
  XOR2_X1 U2984 ( .A(n1581), .B(n1561), .Z(n1582) );
  MUX2_X1 U2985 ( .A(n1603), .B(n1604), .S(n1605), .Z(n1463) );
  XOR2_X1 U2986 ( .A(n1587), .B(n1585), .Z(n1465) );
  XOR2_X1 U2987 ( .A(n1610), .B(n1586), .Z(n1584) );
  XOR2_X1 U2988 ( .A(n1607), .B(n1609), .Z(n1626) );
  XOR2_X1 U2989 ( .A(n1628), .B(n1608), .Z(n1609) );
  XOR2_X1 U2990 ( .A(n1622), .B(n1623), .Z(n1608) );
  XOR2_X1 U2991 ( .A(n1645), .B(n1643), .Z(n1471) );
  XOR2_X1 U2992 ( .A(n1652), .B(n1650), .Z(n1646) );
  XOR2_X1 U2993 ( .A(n1649), .B(n1653), .Z(n1650) );
  MUX2_X1 U2994 ( .A(n1654), .B(n1645), .S(n1655), .Z(n1653) );
  XOR2_X1 U2995 ( .A(n1641), .B(n1642), .Z(n1649) );
  XOR2_X1 U2996 ( .A(n1657), .B(n1635), .Z(n1641) );
  XOR2_X1 U2997 ( .A(n1639), .B(n1634), .Z(n1657) );
  XOR2_X1 U2998 ( .A(n1637), .B(n1659), .Z(n1634) );
  XOR2_X1 U2999 ( .A(n1651), .B(n1644), .Z(n1652) );
  MUX2_X1 U3000 ( .A(n1667), .B(n1668), .S(n1669), .Z(n1651) );
  MUX2_X1 U3001 ( .A(n1675), .B(n1676), .S(n1677), .Z(n1473) );
  XOR2_X1 U3002 ( .A(n1670), .B(n1671), .Z(n1478) );
  XOR2_X1 U3003 ( .A(n1692), .B(n1675), .Z(n1677) );
  MUX2_X1 U3004 ( .A(n1705), .B(n1706), .S(n1707), .Z(n1479) );
  MUX2_X1 U3005 ( .A(n1708), .B(n1709), .S(n1710), .Z(n1482) );
  MUX2_X1 U3006 ( .A(n1712), .B(n1713), .S(n1714), .Z(n1682) );
  XOR2_X1 U3007 ( .A(n1679), .B(n1681), .Z(n1711) );
  XOR2_X1 U3008 ( .A(n1715), .B(n1680), .Z(n1681) );
  XOR2_X1 U3009 ( .A(n1689), .B(n1688), .Z(n1680) );
  XOR2_X1 U3010 ( .A(n1717), .B(n1704), .Z(n1689) );
  XOR2_X1 U3011 ( .A(n1690), .B(n1703), .Z(n1717) );
  XOR2_X1 U3012 ( .A(n1701), .B(n1719), .Z(n1703) );
  MUX2_X1 U3013 ( .A(n1724), .B(n1725), .S(n1726), .Z(n1679) );
  XOR2_X1 U3014 ( .A(n1728), .B(n1710), .Z(n1707) );
  XOR2_X1 U3015 ( .A(n1708), .B(n1729), .Z(n1710) );
  MUX2_X1 U3016 ( .A(n1730), .B(n1731), .S(n1732), .Z(n1729) );
  XOR2_X1 U3017 ( .A(n1712), .B(n1734), .Z(n1714) );
  XOR2_X1 U3018 ( .A(n1726), .B(n1725), .Z(n1734) );
  MUX2_X1 U3019 ( .A(n1741), .B(n1742), .S(n1743), .Z(n1709) );
  MUX2_X1 U3020 ( .A(n1744), .B(n3758), .S(n1745), .Z(n1486) );
  MUX2_X1 U3021 ( .A(n1746), .B(n1747), .S(n1748), .Z(n1485) );
  MUX2_X1 U3022 ( .A(n1749), .B(n1750), .S(n1751), .Z(n1487) );
  MUX2_X1 U3023 ( .A(n1752), .B(n1753), .S(n1754), .Z(n1490) );
  MUX2_X1 U3027 ( .A(n3694), .B(n1773), .S(n1774), .Z(n1491) );
  MUX2_X1 U3028 ( .A(n1775), .B(n1776), .S(n1777), .Z(n1494) );
  XOR2_X1 U3032 ( .A(n1783), .B(n1784), .Z(n1775) );
  MUX2_X1 U3034 ( .A(n1806), .B(n1807), .S(n1808), .Z(n1497) );
  MUX2_X1 U3035 ( .A(n1809), .B(n3719), .S(n1811), .Z(n1499) );
  MUX2_X1 U3036 ( .A(n1812), .B(n1813), .S(n1814), .Z(n1502) );
  XOR2_X1 U3041 ( .A(n1814), .B(n1829), .Z(n1811) );
  XOR2_X1 U3042 ( .A(n1843), .B(n1837), .Z(n1512) );
  XOR2_X1 U3043 ( .A(n1514), .B(n1513), .Z(n1517) );
  XOR2_X1 U3044 ( .A(n1892), .B(n1893), .Z(n1890) );
  XOR2_X1 U3045 ( .A(n1899), .B(n1900), .Z(n1897) );
  XOR2_X1 U3046 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR2_X1 U3047 ( .A(n1907), .B(n1908), .Z(n1906) );
  XOR2_X1 U3048 ( .A(n1911), .B(n1912), .Z(n1910) );
  XOR2_X1 U3049 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR2_X1 U3050 ( .A(n1919), .B(n1920), .Z(n1918) );
  XOR2_X1 U3051 ( .A(n1923), .B(n1924), .Z(n1922) );
  XOR2_X1 U3052 ( .A(n1925), .B(n1926), .Z(p6_S[45]) );
  XOR2_X1 U3054 ( .A(n1935), .B(n1936), .Z(n1934) );
  XOR2_X1 U3060 ( .A(n1957), .B(n1958), .Z(n1956) );
  XOR2_X1 U3061 ( .A(n3710), .B(n1960), .Z(p6_S[36]) );
  XOR2_X1 U3062 ( .A(n1961), .B(n1962), .Z(n1960) );
  XOR2_X1 U3064 ( .A(n3711), .B(n1974), .Z(n1971) );
  XOR2_X1 U3065 ( .A(n1975), .B(n1976), .Z(p6_S[33]) );
  XOR2_X1 U3067 ( .A(n3757), .B(n1987), .Z(n1898) );
  XOR2_X1 U3068 ( .A(n1986), .B(n1985), .Z(n1987) );
  XOR2_X1 U3069 ( .A(n2002), .B(n1992), .Z(n2000) );
  MUX2_X1 U3070 ( .A(n2013), .B(n2014), .S(n2015), .Z(n1903) );
  XOR2_X1 U3071 ( .A(n2011), .B(n2009), .Z(n1905) );
  XOR2_X1 U3072 ( .A(n2016), .B(n2010), .Z(n2009) );
  MUX2_X1 U3073 ( .A(n2038), .B(n2039), .S(n2040), .Z(n1912) );
  XOR2_X1 U3074 ( .A(n2028), .B(n2026), .Z(n1911) );
  XOR2_X1 U3075 ( .A(n2043), .B(n2027), .Z(n2025) );
  XOR2_X1 U3076 ( .A(n2032), .B(n2033), .Z(n2043) );
  XOR2_X1 U3077 ( .A(n2031), .B(n2011), .Z(n2032) );
  MUX2_X1 U3078 ( .A(n2053), .B(n2054), .S(n2055), .Z(n1913) );
  XOR2_X1 U3079 ( .A(n2037), .B(n2035), .Z(n1915) );
  XOR2_X1 U3080 ( .A(n2060), .B(n2036), .Z(n2034) );
  XOR2_X1 U3081 ( .A(n2057), .B(n2059), .Z(n2076) );
  XOR2_X1 U3082 ( .A(n2078), .B(n2058), .Z(n2059) );
  XOR2_X1 U3083 ( .A(n2072), .B(n2073), .Z(n2058) );
  XOR2_X1 U3084 ( .A(n2095), .B(n2093), .Z(n1921) );
  XOR2_X1 U3085 ( .A(n2102), .B(n2100), .Z(n2096) );
  XOR2_X1 U3086 ( .A(n2099), .B(n2103), .Z(n2100) );
  MUX2_X1 U3087 ( .A(n2104), .B(n2095), .S(n2105), .Z(n2103) );
  XOR2_X1 U3088 ( .A(n2091), .B(n2092), .Z(n2099) );
  XOR2_X1 U3089 ( .A(n2107), .B(n2085), .Z(n2091) );
  XOR2_X1 U3090 ( .A(n2089), .B(n2084), .Z(n2107) );
  XOR2_X1 U3091 ( .A(n2087), .B(n2109), .Z(n2084) );
  XOR2_X1 U3092 ( .A(n2101), .B(n2094), .Z(n2102) );
  MUX2_X1 U3093 ( .A(n2117), .B(n2118), .S(n2119), .Z(n2101) );
  MUX2_X1 U3094 ( .A(n2125), .B(n2126), .S(n2127), .Z(n1923) );
  XOR2_X1 U3095 ( .A(n2120), .B(n2121), .Z(n1928) );
  XOR2_X1 U3096 ( .A(n2142), .B(n2125), .Z(n2127) );
  MUX2_X1 U3097 ( .A(n2155), .B(n2156), .S(n2157), .Z(n1929) );
  MUX2_X1 U3098 ( .A(n2158), .B(n2159), .S(n2160), .Z(n1932) );
  MUX2_X1 U3099 ( .A(n2162), .B(n2163), .S(n2164), .Z(n2132) );
  XOR2_X1 U3102 ( .A(n2139), .B(n2138), .Z(n2130) );
  XOR2_X1 U3103 ( .A(n2167), .B(n2154), .Z(n2139) );
  XOR2_X1 U3104 ( .A(n2140), .B(n2153), .Z(n2167) );
  XOR2_X1 U3105 ( .A(n2151), .B(n2169), .Z(n2153) );
  MUX2_X1 U3106 ( .A(n2174), .B(n2175), .S(n2176), .Z(n2129) );
  XOR2_X1 U3107 ( .A(n2178), .B(n2160), .Z(n2157) );
  XOR2_X1 U3108 ( .A(n2158), .B(n2179), .Z(n2160) );
  MUX2_X1 U3109 ( .A(n2180), .B(n2181), .S(n2182), .Z(n2179) );
  XOR2_X1 U3110 ( .A(n2162), .B(n2184), .Z(n2164) );
  XOR2_X1 U3111 ( .A(n2176), .B(n2175), .Z(n2184) );
  MUX2_X1 U3112 ( .A(n2191), .B(n2192), .S(n2193), .Z(n2159) );
  MUX2_X1 U3113 ( .A(n2194), .B(n3757), .S(n2195), .Z(n1936) );
  MUX2_X1 U3114 ( .A(n2196), .B(n2197), .S(n2198), .Z(n1935) );
  MUX2_X1 U3115 ( .A(n2199), .B(n2200), .S(n2201), .Z(n1937) );
  MUX2_X1 U3116 ( .A(n2202), .B(n2203), .S(n2204), .Z(n1940) );
  MUX2_X1 U3120 ( .A(n3674), .B(n2223), .S(n2224), .Z(n1941) );
  MUX2_X1 U3121 ( .A(n2225), .B(n2226), .S(n2227), .Z(n1944) );
  XOR2_X1 U3124 ( .A(n2247), .B(n2225), .Z(n2227) );
  XOR2_X1 U3125 ( .A(n2233), .B(n2234), .Z(n2225) );
  MUX2_X1 U3126 ( .A(n2253), .B(n2254), .S(n2255), .Z(n1948) );
  MUX2_X1 U3127 ( .A(n2256), .B(n2257), .S(n2258), .Z(n1947) );
  MUX2_X1 U3128 ( .A(n2259), .B(n3713), .S(n2261), .Z(n1949) );
  MUX2_X1 U3129 ( .A(n2262), .B(n2263), .S(n2264), .Z(n1952) );
  XOR2_X1 U3135 ( .A(n2293), .B(n2287), .Z(n1962) );
  XOR2_X1 U3137 ( .A(n2342), .B(n2343), .Z(n2340) );
  XOR2_X1 U3138 ( .A(n2349), .B(n2350), .Z(n2347) );
  XOR2_X1 U3139 ( .A(n2353), .B(n2354), .Z(n2352) );
  XOR2_X1 U3140 ( .A(n2357), .B(n2358), .Z(n2356) );
  XOR2_X1 U3141 ( .A(n2361), .B(n2362), .Z(n2360) );
  XOR2_X1 U3142 ( .A(n2365), .B(n2366), .Z(n2364) );
  XOR2_X1 U3143 ( .A(n2369), .B(n2370), .Z(n2368) );
  XOR2_X1 U3144 ( .A(n2373), .B(n2374), .Z(n2372) );
  XOR2_X1 U3145 ( .A(n2375), .B(n2376), .Z(p11_S[45]) );
  XOR2_X1 U3149 ( .A(n2393), .B(n2394), .Z(n2392) );
  XOR2_X1 U3150 ( .A(n2397), .B(n2398), .Z(n2396) );
  XOR2_X1 U3151 ( .A(n2401), .B(n2402), .Z(n2400) );
  XOR2_X1 U3152 ( .A(n2403), .B(n2404), .Z(p11_S[38]) );
  XOR2_X1 U3153 ( .A(n2405), .B(n2406), .Z(p11_S[37]) );
  XOR2_X1 U3154 ( .A(n2407), .B(n2408), .Z(n2406) );
  XOR2_X1 U3155 ( .A(n2415), .B(n2416), .Z(p11_S[35]) );
  XOR2_X1 U3156 ( .A(n2423), .B(n2424), .Z(n2421) );
  XOR2_X1 U3157 ( .A(n2425), .B(n2426), .Z(p11_S[33]) );
  XOR2_X1 U3159 ( .A(n2444), .B(n2437), .Z(n2348) );
  XOR2_X1 U3160 ( .A(n2436), .B(n2435), .Z(n2437) );
  XOR2_X1 U3161 ( .A(n2452), .B(n2442), .Z(n2450) );
  MUX2_X1 U3162 ( .A(n2463), .B(n2464), .S(n2465), .Z(n2353) );
  XOR2_X1 U3163 ( .A(n2461), .B(n2459), .Z(n2355) );
  XOR2_X1 U3164 ( .A(n2466), .B(n2460), .Z(n2459) );
  MUX2_X1 U3165 ( .A(n2488), .B(n2489), .S(n2490), .Z(n2362) );
  XOR2_X1 U3166 ( .A(n2478), .B(n2476), .Z(n2361) );
  XOR2_X1 U3167 ( .A(n2493), .B(n2477), .Z(n2475) );
  XOR2_X1 U3168 ( .A(n2482), .B(n2483), .Z(n2493) );
  XOR2_X1 U3169 ( .A(n2481), .B(n2461), .Z(n2482) );
  MUX2_X1 U3170 ( .A(n2503), .B(n2504), .S(n2505), .Z(n2363) );
  XOR2_X1 U3171 ( .A(n2487), .B(n2485), .Z(n2365) );
  XOR2_X1 U3172 ( .A(n2510), .B(n2486), .Z(n2484) );
  XOR2_X1 U3173 ( .A(n2507), .B(n2509), .Z(n2526) );
  XOR2_X1 U3174 ( .A(n2528), .B(n2508), .Z(n2509) );
  XOR2_X1 U3175 ( .A(n2522), .B(n2523), .Z(n2508) );
  XOR2_X1 U3176 ( .A(n2545), .B(n2543), .Z(n2371) );
  XOR2_X1 U3177 ( .A(n2552), .B(n2550), .Z(n2546) );
  MUX2_X1 U3179 ( .A(n2554), .B(n2545), .S(n2555), .Z(n2553) );
  XOR2_X1 U3180 ( .A(n2541), .B(n2542), .Z(n2549) );
  XOR2_X1 U3181 ( .A(n2557), .B(n2535), .Z(n2541) );
  XOR2_X1 U3182 ( .A(n2539), .B(n2534), .Z(n2557) );
  XOR2_X1 U3183 ( .A(n2537), .B(n2559), .Z(n2534) );
  XOR2_X1 U3184 ( .A(n2551), .B(n2544), .Z(n2552) );
  MUX2_X1 U3185 ( .A(n2567), .B(n2568), .S(n2569), .Z(n2551) );
  MUX2_X1 U3186 ( .A(n2575), .B(n2576), .S(n2577), .Z(n2373) );
  XOR2_X1 U3187 ( .A(n2570), .B(n2571), .Z(n2377) );
  XOR2_X1 U3188 ( .A(n2575), .B(n2592), .Z(n2577) );
  MUX2_X1 U3189 ( .A(n2593), .B(n2594), .S(n2595), .Z(n2592) );
  MUX2_X1 U3190 ( .A(n2604), .B(n2605), .S(n2606), .Z(n2379) );
  MUX2_X1 U3191 ( .A(n2607), .B(n2608), .S(n2609), .Z(n2382) );
  XOR2_X1 U3194 ( .A(n2581), .B(n2582), .Z(n2610) );
  XOR2_X1 U3196 ( .A(n2590), .B(n2589), .Z(n2580) );
  XOR2_X1 U3197 ( .A(n2621), .B(n2593), .Z(n2590) );
  XOR2_X1 U3198 ( .A(n2588), .B(n2595), .Z(n2621) );
  XOR2_X1 U3199 ( .A(n2594), .B(n2623), .Z(n2595) );
  XOR2_X1 U3200 ( .A(n2631), .B(n2605), .Z(n2606) );
  XOR2_X1 U3201 ( .A(n2607), .B(n2633), .Z(n2609) );
  MUX2_X1 U3202 ( .A(n2634), .B(n2635), .S(n2636), .Z(n2633) );
  XOR2_X1 U3203 ( .A(n2614), .B(n2613), .Z(n2607) );
  MUX2_X1 U3204 ( .A(n2644), .B(n2645), .S(n2646), .Z(n2608) );
  MUX2_X1 U3205 ( .A(n2647), .B(n2444), .S(n2648), .Z(n2386) );
  MUX2_X1 U3206 ( .A(n2649), .B(n2650), .S(n2651), .Z(n2385) );
  MUX2_X1 U3207 ( .A(n2652), .B(n2653), .S(n2654), .Z(n2387) );
  MUX2_X1 U3208 ( .A(n2655), .B(n2656), .S(n2657), .Z(n2390) );
  XOR2_X1 U3211 ( .A(n2646), .B(n2645), .Z(n2650) );
  MUX2_X1 U3212 ( .A(n2674), .B(n2675), .S(n2676), .Z(n2391) );
  MUX2_X1 U3213 ( .A(n2677), .B(n2678), .S(n2679), .Z(n2394) );
  XOR2_X1 U3214 ( .A(n2654), .B(n2653), .Z(n2393) );
  XOR2_X1 U3217 ( .A(n2685), .B(n2686), .Z(n2677) );
  MUX2_X1 U3218 ( .A(n2705), .B(n2706), .S(n2707), .Z(n2398) );
  MUX2_X1 U3219 ( .A(n2708), .B(n2709), .S(n2710), .Z(n2397) );
  MUX2_X1 U3220 ( .A(n2711), .B(n2712), .S(n2713), .Z(n2399) );
  MUX2_X1 U3221 ( .A(n2714), .B(n2715), .S(n2716), .Z(n2402) );
  XOR2_X1 U3222 ( .A(n2707), .B(n2706), .Z(n2401) );
  XOR2_X1 U3223 ( .A(n2705), .B(n2718), .Z(n2707) );
  XOR2_X1 U3224 ( .A(n2709), .B(n2710), .Z(n2718) );
  XOR2_X1 U3225 ( .A(n2719), .B(n2708), .Z(n2710) );
  XOR2_X1 U3227 ( .A(n2414), .B(n2413), .Z(n2417) );
  XOR2_X1 U3228 ( .A(n2792), .B(n2793), .Z(n2790) );
  XOR2_X1 U3229 ( .A(n2799), .B(n2800), .Z(n2797) );
  XOR2_X1 U3230 ( .A(n2803), .B(n2804), .Z(n2802) );
  XOR2_X1 U3231 ( .A(n2807), .B(n2808), .Z(n2806) );
  XOR2_X1 U3232 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR2_X1 U3233 ( .A(n2815), .B(n2816), .Z(n2814) );
  XOR2_X1 U3234 ( .A(n2819), .B(n2820), .Z(n2818) );
  XOR2_X1 U3235 ( .A(n2823), .B(n2824), .Z(n2822) );
  XOR2_X1 U3236 ( .A(n2825), .B(n2826), .Z(p10_S[45]) );
  XOR2_X1 U3238 ( .A(n2835), .B(n2836), .Z(n2834) );
  XOR2_X1 U3240 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR2_X1 U3242 ( .A(n2851), .B(n2852), .Z(n2850) );
  XOR2_X1 U3243 ( .A(n2853), .B(n2854), .Z(p10_S[38]) );
  XOR2_X1 U3244 ( .A(n2855), .B(n2856), .Z(p10_S[37]) );
  XOR2_X1 U3245 ( .A(n2857), .B(n2858), .Z(n2856) );
  XOR2_X1 U3246 ( .A(n2865), .B(n2866), .Z(p10_S[35]) );
  XOR2_X1 U3247 ( .A(n2873), .B(n2874), .Z(n2871) );
  XOR2_X1 U3248 ( .A(n2875), .B(n2876), .Z(p10_S[33]) );
  XOR2_X1 U3250 ( .A(n2894), .B(n2887), .Z(n2798) );
  XOR2_X1 U3251 ( .A(n2886), .B(n2885), .Z(n2887) );
  XOR2_X1 U3252 ( .A(n2902), .B(n2892), .Z(n2900) );
  MUX2_X1 U3253 ( .A(n2913), .B(n2914), .S(n2915), .Z(n2803) );
  XOR2_X1 U3254 ( .A(n2911), .B(n2909), .Z(n2805) );
  XOR2_X1 U3255 ( .A(n2916), .B(n2910), .Z(n2909) );
  MUX2_X1 U3256 ( .A(n2938), .B(n2939), .S(n2940), .Z(n2812) );
  XOR2_X1 U3257 ( .A(n2928), .B(n2926), .Z(n2811) );
  XOR2_X1 U3258 ( .A(n2943), .B(n2927), .Z(n2925) );
  XOR2_X1 U3259 ( .A(n2932), .B(n2933), .Z(n2943) );
  XOR2_X1 U3260 ( .A(n2931), .B(n2911), .Z(n2932) );
  MUX2_X1 U3261 ( .A(n2953), .B(n2954), .S(n2955), .Z(n2813) );
  XOR2_X1 U3262 ( .A(n2937), .B(n2935), .Z(n2815) );
  XOR2_X1 U3263 ( .A(n2960), .B(n2936), .Z(n2934) );
  XOR2_X1 U3264 ( .A(n2957), .B(n2959), .Z(n2976) );
  XOR2_X1 U3265 ( .A(n2958), .B(n2978), .Z(n2959) );
  MUX2_X1 U3266 ( .A(n2979), .B(n2980), .S(n2981), .Z(n2978) );
  XOR2_X1 U3267 ( .A(n2972), .B(n2973), .Z(n2958) );
  XOR2_X1 U3268 ( .A(n2994), .B(n2992), .Z(n2821) );
  XOR2_X1 U3269 ( .A(n3001), .B(n2999), .Z(n2995) );
  XOR2_X1 U3270 ( .A(n2998), .B(n3002), .Z(n2999) );
  MUX2_X1 U3271 ( .A(n3003), .B(n2994), .S(n3004), .Z(n3002) );
  XOR2_X1 U3272 ( .A(n2990), .B(n2991), .Z(n2998) );
  XOR2_X1 U3273 ( .A(n3006), .B(n2981), .Z(n2990) );
  XOR2_X1 U3274 ( .A(n3000), .B(n2993), .Z(n3001) );
  MUX2_X1 U3275 ( .A(n3016), .B(n3017), .S(n3018), .Z(n3000) );
  MUX2_X1 U3276 ( .A(n3024), .B(n3025), .S(n3026), .Z(n2823) );
  XOR2_X1 U3277 ( .A(n3019), .B(n3020), .Z(n2828) );
  XOR2_X1 U3278 ( .A(n3024), .B(n3040), .Z(n3026) );
  MUX2_X1 U3279 ( .A(n3041), .B(n3042), .S(n3043), .Z(n3040) );
  MUX2_X1 U3281 ( .A(n3055), .B(n3056), .S(n3057), .Z(n2832) );
  MUX2_X1 U3282 ( .A(n3059), .B(n3060), .S(n3061), .Z(n3031) );
  XOR2_X1 U3283 ( .A(n3028), .B(n3030), .Z(n3058) );
  XOR2_X1 U3284 ( .A(n3062), .B(n3029), .Z(n3030) );
  XOR2_X1 U3285 ( .A(n3038), .B(n3037), .Z(n3029) );
  XOR2_X1 U3286 ( .A(n3064), .B(n3041), .Z(n3038) );
  XOR2_X1 U3287 ( .A(n3036), .B(n3043), .Z(n3064) );
  XOR2_X1 U3288 ( .A(n3042), .B(n3066), .Z(n3043) );
  MUX2_X1 U3289 ( .A(n3073), .B(n3074), .S(n3075), .Z(n3028) );
  XOR2_X1 U3290 ( .A(n3077), .B(n3053), .Z(n3054) );
  XOR2_X1 U3291 ( .A(n3055), .B(n3079), .Z(n3057) );
  MUX2_X1 U3292 ( .A(n3080), .B(n3081), .S(n3082), .Z(n3079) );
  XOR2_X1 U3293 ( .A(n3059), .B(n3084), .Z(n3061) );
  XOR2_X1 U3294 ( .A(n3075), .B(n3074), .Z(n3084) );
  MUX2_X1 U3295 ( .A(n3090), .B(n3091), .S(n3092), .Z(n3056) );
  MUX2_X1 U3296 ( .A(n3093), .B(n2894), .S(n3094), .Z(n2836) );
  MUX2_X1 U3297 ( .A(n3095), .B(n3096), .S(n3097), .Z(n2835) );
  MUX2_X1 U3298 ( .A(n3098), .B(n3099), .S(n3100), .Z(n2837) );
  MUX2_X1 U3299 ( .A(n3101), .B(n3102), .S(n3103), .Z(n2840) );
  XOR2_X1 U3302 ( .A(n3092), .B(n3091), .Z(n3096) );
  MUX2_X1 U3303 ( .A(n3120), .B(n3121), .S(n3122), .Z(n2841) );
  MUX2_X1 U3304 ( .A(n3123), .B(n3124), .S(n3125), .Z(n2844) );
  XOR2_X1 U3305 ( .A(n3100), .B(n3099), .Z(n2843) );
  XOR2_X1 U3308 ( .A(n3131), .B(n3132), .Z(n3123) );
  MUX2_X1 U3310 ( .A(n3154), .B(n3155), .S(n3156), .Z(n2847) );
  MUX2_X1 U3311 ( .A(n3157), .B(n3158), .S(n3159), .Z(n2849) );
  MUX2_X1 U3312 ( .A(n3160), .B(n3161), .S(n3162), .Z(n2852) );
  XOR2_X1 U3313 ( .A(n3153), .B(n3152), .Z(n2851) );
  XOR2_X1 U3316 ( .A(n3165), .B(n3154), .Z(n3156) );
  XOR2_X1 U3317 ( .A(n3162), .B(n3177), .Z(n3159) );
  MUX2_X1 U3320 ( .A(DIN[13]), .B(xin_in[13]), .S(n3850), .Z(n45) );
  MUX2_X1 U3321 ( .A(DIN[12]), .B(xin_in[12]), .S(n3846), .Z(n44) );
  MUX2_X1 U3322 ( .A(DIN[11]), .B(xin_in[11]), .S(n3852), .Z(n43) );
  MUX2_X1 U3323 ( .A(DIN[10]), .B(xin_in[10]), .S(n3850), .Z(n42) );
  MUX2_X1 U3324 ( .A(DIN[9]), .B(xin_in[9]), .S(n3848), .Z(n41) );
  MUX2_X1 U3325 ( .A(DIN[8]), .B(xin_in[8]), .S(n3852), .Z(n40) );
  MUX2_X1 U3326 ( .A(DIN[7]), .B(xin_in[7]), .S(n3848), .Z(n39) );
  MUX2_X1 U3327 ( .A(DIN[6]), .B(xin_in[6]), .S(n3848), .Z(n38) );
  MUX2_X1 U3328 ( .A(DIN[5]), .B(xin_in[5]), .S(n3849), .Z(n37) );
  MUX2_X1 U3329 ( .A(DIN[4]), .B(xin_in[4]), .S(n3851), .Z(n36) );
  MUX2_X1 U3330 ( .A(DIN[3]), .B(xin_in[3]), .S(n3847), .Z(n35) );
  MUX2_X1 U3331 ( .A(DIN[2]), .B(xin_in[2]), .S(n3852), .Z(n34) );
  MUX2_X1 U3332 ( .A(DIN[1]), .B(xin_in[1]), .S(n3847), .Z(n33) );
  MUX2_X1 U3333 ( .A(DIN[0]), .B(xin_in[0]), .S(n3847), .Z(n32) );
  XOR2_X1 U3334 ( .A(reg7[12]), .B(n3241), .Z(SUB1_N12) );
  XOR2_X1 U3335 ( .A(n3748), .B(n3242), .Z(SUB1_N11) );
  MUX2_X1 U3336 ( .A(xin_in[13]), .B(xin[13]), .S(n3849), .Z(REGISTER_in_n42)
         );
  MUX2_X1 U3337 ( .A(xin_in[12]), .B(xin[12]), .S(n3851), .Z(REGISTER_in_n41)
         );
  MUX2_X1 U3338 ( .A(xin_in[11]), .B(xin[11]), .S(n3847), .Z(REGISTER_in_n40)
         );
  MUX2_X1 U3339 ( .A(xin_in[10]), .B(xin[10]), .S(n3848), .Z(REGISTER_in_n39)
         );
  MUX2_X1 U3340 ( .A(xin_in[9]), .B(xin[9]), .S(n3848), .Z(REGISTER_in_n38) );
  MUX2_X1 U3341 ( .A(xin_in[8]), .B(xin[8]), .S(n3849), .Z(REGISTER_in_n37) );
  MUX2_X1 U3342 ( .A(xin_in[7]), .B(xin[7]), .S(n3849), .Z(REGISTER_in_n36) );
  MUX2_X1 U3343 ( .A(xin_in[6]), .B(xin[6]), .S(n3852), .Z(REGISTER_in_n35) );
  MUX2_X1 U3344 ( .A(xin_in[5]), .B(xin[5]), .S(n3847), .Z(REGISTER_in_n34) );
  MUX2_X1 U3345 ( .A(xin_in[4]), .B(xin[4]), .S(n3850), .Z(REGISTER_in_n33) );
  MUX2_X1 U3346 ( .A(xin_in[3]), .B(xin[3]), .S(n3846), .Z(REGISTER_in_n32) );
  MUX2_X1 U3347 ( .A(xin_in[2]), .B(xin[2]), .S(n3851), .Z(REGISTER_in_n31) );
  MUX2_X1 U3348 ( .A(xin_in[1]), .B(xin[1]), .S(n3850), .Z(REGISTER_in_n30) );
  MUX2_X1 U3349 ( .A(xin_in[0]), .B(xin[0]), .S(n3849), .Z(REGISTER_in_n29) );
  MUX2_X1 U3350 ( .A(temp6[0]), .B(reg7[0]), .S(n3851), .Z(REG61_n62) );
  MUX2_X1 U3351 ( .A(temp6[1]), .B(reg7[1]), .S(n3846), .Z(REG61_n61) );
  MUX2_X1 U3352 ( .A(temp6[2]), .B(reg7[2]), .S(n3850), .Z(REG61_n60) );
  MUX2_X1 U3353 ( .A(temp6[3]), .B(reg7[3]), .S(n3849), .Z(REG61_n59) );
  MUX2_X1 U3355 ( .A(temp6[5]), .B(reg7[5]), .S(n3852), .Z(REG61_n57) );
  MUX2_X1 U3356 ( .A(temp6[6]), .B(reg7[6]), .S(n3847), .Z(REG61_n56) );
  MUX2_X1 U3357 ( .A(temp6[7]), .B(reg7[7]), .S(n3852), .Z(REG61_n55) );
  MUX2_X1 U3358 ( .A(temp6[8]), .B(reg7[8]), .S(n3850), .Z(REG61_n54) );
  MUX2_X1 U3359 ( .A(temp6[9]), .B(reg7[9]), .S(n3846), .Z(REG61_n53) );
  MUX2_X1 U3360 ( .A(temp6[10]), .B(reg7[10]), .S(n3848), .Z(REG61_n52) );
  MUX2_X1 U3361 ( .A(temp6[11]), .B(reg7[11]), .S(n3846), .Z(REG61_n51) );
  MUX2_X1 U3362 ( .A(temp6[12]), .B(reg7[12]), .S(n3851), .Z(REG61_n50) );
  MUX2_X1 U3364 ( .A(temp5[0]), .B(reg6[0]), .S(n3846), .Z(REG51_n63) );
  MUX2_X1 U3365 ( .A(temp5[1]), .B(reg6[1]), .S(n3852), .Z(REG51_n62) );
  MUX2_X1 U3366 ( .A(temp5[2]), .B(reg6[2]), .S(n3850), .Z(REG51_n61) );
  MUX2_X1 U3367 ( .A(temp5[3]), .B(reg6[3]), .S(n3852), .Z(REG51_n60) );
  MUX2_X1 U3368 ( .A(temp5[4]), .B(reg6[4]), .S(n3850), .Z(REG51_n59) );
  MUX2_X1 U3369 ( .A(temp5[5]), .B(reg6[5]), .S(n3849), .Z(REG51_n58) );
  MUX2_X1 U3370 ( .A(temp5[6]), .B(reg6[6]), .S(n3852), .Z(REG51_n57) );
  MUX2_X1 U3371 ( .A(temp5[7]), .B(reg6[7]), .S(n3850), .Z(REG51_n56) );
  MUX2_X1 U3372 ( .A(temp5[8]), .B(reg6[8]), .S(n3848), .Z(REG51_n55) );
  MUX2_X1 U3373 ( .A(temp5[9]), .B(reg6[9]), .S(n3850), .Z(REG51_n54) );
  MUX2_X1 U3374 ( .A(temp5[10]), .B(reg6[10]), .S(n3849), .Z(REG51_n53) );
  MUX2_X1 U3375 ( .A(temp5[11]), .B(reg6[11]), .S(n3846), .Z(REG51_n52) );
  MUX2_X1 U3376 ( .A(temp5[12]), .B(reg6[12]), .S(n3846), .Z(REG51_n51) );
  MUX2_X1 U3378 ( .A(temp4[0]), .B(mul4_reg[0]), .S(n3848), .Z(REG4_1_n62) );
  MUX2_X1 U3379 ( .A(temp4[1]), .B(mul4_reg[1]), .S(n3849), .Z(REG4_1_n61) );
  MUX2_X1 U3380 ( .A(temp4[2]), .B(mul4_reg[2]), .S(n3851), .Z(REG4_1_n60) );
  MUX2_X1 U3381 ( .A(temp4[3]), .B(mul4_reg[3]), .S(n3850), .Z(REG4_1_n59) );
  MUX2_X1 U3382 ( .A(temp4[4]), .B(mul4_reg[4]), .S(n3847), .Z(REG4_1_n58) );
  MUX2_X1 U3383 ( .A(temp4[5]), .B(mul4_reg[5]), .S(n3851), .Z(REG4_1_n57) );
  MUX2_X1 U3384 ( .A(temp4[6]), .B(mul4_reg[6]), .S(n3847), .Z(REG4_1_n56) );
  MUX2_X1 U3385 ( .A(temp4[7]), .B(mul4_reg[7]), .S(n3851), .Z(REG4_1_n55) );
  MUX2_X1 U3386 ( .A(temp4[8]), .B(mul4_reg[8]), .S(n3852), .Z(REG4_1_n54) );
  MUX2_X1 U3387 ( .A(temp4[9]), .B(mul4_reg[9]), .S(n3849), .Z(REG4_1_n53) );
  MUX2_X1 U3388 ( .A(temp4[10]), .B(mul4_reg[10]), .S(n3851), .Z(REG4_1_n52)
         );
  MUX2_X1 U3389 ( .A(temp4[11]), .B(mul4_reg[11]), .S(n3852), .Z(REG4_1_n51)
         );
  MUX2_X1 U3392 ( .A(temp3[0]), .B(mul3_reg[0]), .S(n3847), .Z(REG3_1_n62) );
  MUX2_X1 U3393 ( .A(temp3[1]), .B(mul3_reg[1]), .S(n3851), .Z(REG3_1_n61) );
  MUX2_X1 U3394 ( .A(temp3[2]), .B(mul3_reg[2]), .S(n3850), .Z(REG3_1_n60) );
  MUX2_X1 U3395 ( .A(temp3[3]), .B(mul3_reg[3]), .S(n3852), .Z(REG3_1_n59) );
  MUX2_X1 U3396 ( .A(temp3[4]), .B(mul3_reg[4]), .S(n3849), .Z(REG3_1_n58) );
  MUX2_X1 U3397 ( .A(temp3[5]), .B(mul3_reg[5]), .S(n3847), .Z(REG3_1_n57) );
  MUX2_X1 U3398 ( .A(temp3[6]), .B(mul3_reg[6]), .S(n3850), .Z(REG3_1_n56) );
  MUX2_X1 U3399 ( .A(temp3[7]), .B(mul3_reg[7]), .S(n3849), .Z(REG3_1_n55) );
  MUX2_X1 U3400 ( .A(temp3[8]), .B(mul3_reg[8]), .S(n3848), .Z(REG3_1_n54) );
  MUX2_X1 U3401 ( .A(temp3[9]), .B(mul3_reg[9]), .S(n3850), .Z(REG3_1_n53) );
  MUX2_X1 U3402 ( .A(temp3[10]), .B(mul3_reg[10]), .S(n3846), .Z(REG3_1_n52)
         );
  MUX2_X1 U3403 ( .A(temp3[11]), .B(mul3_reg[11]), .S(n3851), .Z(REG3_1_n51)
         );
  MUX2_X1 U3406 ( .A(temp2[0]), .B(mul2_reg[0]), .S(n3851), .Z(REG2_1_n62) );
  MUX2_X1 U3407 ( .A(temp2[1]), .B(mul2_reg[1]), .S(n3848), .Z(REG2_1_n61) );
  MUX2_X1 U3408 ( .A(temp2[2]), .B(mul2_reg[2]), .S(n3849), .Z(REG2_1_n60) );
  MUX2_X1 U3409 ( .A(temp2[3]), .B(mul2_reg[3]), .S(n3847), .Z(REG2_1_n59) );
  MUX2_X1 U3410 ( .A(temp2[4]), .B(mul2_reg[4]), .S(n3847), .Z(REG2_1_n58) );
  MUX2_X1 U3411 ( .A(temp2[5]), .B(mul2_reg[5]), .S(n3852), .Z(REG2_1_n57) );
  MUX2_X1 U3412 ( .A(temp2[6]), .B(mul2_reg[6]), .S(n3848), .Z(REG2_1_n56) );
  MUX2_X1 U3413 ( .A(temp2[7]), .B(mul2_reg[7]), .S(n3846), .Z(REG2_1_n55) );
  MUX2_X1 U3414 ( .A(temp2[8]), .B(mul2_reg[8]), .S(n3846), .Z(REG2_1_n54) );
  MUX2_X1 U3415 ( .A(temp2[9]), .B(mul2_reg[9]), .S(n3846), .Z(REG2_1_n53) );
  MUX2_X1 U3416 ( .A(temp2[10]), .B(mul2_reg[10]), .S(n3847), .Z(REG2_1_n52)
         );
  MUX2_X1 U3417 ( .A(temp2[11]), .B(mul2_reg[11]), .S(n3847), .Z(REG2_1_n51)
         );
  MUX2_X1 U3418 ( .A(temp2[12]), .B(mul2_reg[12]), .S(n3847), .Z(REG2_1_n50)
         );
  MUX2_X1 U3420 ( .A(temp1[0]), .B(mul1_reg[0]), .S(n3848), .Z(REG1_1_n62) );
  MUX2_X1 U3421 ( .A(temp1[1]), .B(mul1_reg[1]), .S(n3848), .Z(REG1_1_n61) );
  MUX2_X1 U3422 ( .A(temp1[2]), .B(mul1_reg[2]), .S(n3849), .Z(REG1_1_n60) );
  MUX2_X1 U3423 ( .A(temp1[3]), .B(mul1_reg[3]), .S(n3849), .Z(REG1_1_n59) );
  MUX2_X1 U3424 ( .A(temp1[4]), .B(mul1_reg[4]), .S(n3849), .Z(REG1_1_n58) );
  MUX2_X1 U3425 ( .A(temp1[5]), .B(mul1_reg[5]), .S(n3850), .Z(REG1_1_n57) );
  MUX2_X1 U3426 ( .A(temp1[6]), .B(mul1_reg[6]), .S(n3850), .Z(REG1_1_n56) );
  MUX2_X1 U3427 ( .A(temp1[7]), .B(mul1_reg[7]), .S(n3850), .Z(REG1_1_n55) );
  MUX2_X1 U3428 ( .A(temp1[8]), .B(mul1_reg[8]), .S(n3851), .Z(REG1_1_n54) );
  MUX2_X1 U3429 ( .A(temp1[9]), .B(mul1_reg[9]), .S(n3851), .Z(REG1_1_n53) );
  MUX2_X1 U3430 ( .A(temp1[10]), .B(mul1_reg[10]), .S(n3851), .Z(REG1_1_n52)
         );
  MUX2_X1 U3431 ( .A(temp1[11]), .B(mul1_reg[11]), .S(n3852), .Z(REG1_1_n51)
         );
  MUX2_X1 U3432 ( .A(temp1[12]), .B(mul1_reg[12]), .S(n3852), .Z(REG1_1_n50)
         );
  MUX2_X1 U3363 ( .A(temp6[13]), .B(reg7[13]), .S(n3848), .Z(REG61_n49) );
  MUX2_X1 U3433 ( .A(temp1[13]), .B(mul1_reg[13]), .S(n3852), .Z(REG1_1_n49)
         );
  XOR2_X1 U3055 ( .A(n1939), .B(n1940), .Z(n1938) );
  MUX2_X1 U3377 ( .A(temp5[13]), .B(reg6[13]), .S(n3851), .Z(REG51_n50) );
  MUX2_X1 U3391 ( .A(temp4[13]), .B(mul4_reg[13]), .S(n3852), .Z(REG4_1_n49)
         );
  XOR2_X1 U2776 ( .A(n590), .B(n591), .Z(n589) );
  XOR2_X1 U2778 ( .A(n598), .B(n599), .Z(n597) );
  MUX2_X1 U3405 ( .A(temp3[13]), .B(mul3_reg[13]), .S(n3846), .Z(REG3_1_n49)
         );
  XOR2_X1 U3241 ( .A(n2847), .B(n2848), .Z(n2846) );
  MUX2_X1 U3309 ( .A(n3151), .B(n3152), .S(n3153), .Z(n2848) );
  XOR2_X1 U2872 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR2_X1 U2944 ( .A(n1355), .B(n1354), .Z(n1052) );
  XOR2_X1 U2869 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR2_X1 U3300 ( .A(n3097), .B(n3093), .Z(n3105) );
  MUX2_X1 U3419 ( .A(temp2[13]), .B(mul2_reg[13]), .S(n3848), .Z(REG2_1_n49)
         );
  XOR2_X1 U2964 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR2_X1 U3057 ( .A(n1947), .B(n1948), .Z(n1946) );
  XOR2_X1 U2931 ( .A(n1299), .B(n1295), .Z(n1307) );
  XOR2_X1 U2839 ( .A(n862), .B(n848), .Z(n849) );
  XOR2_X1 U3118 ( .A(n2211), .B(n2197), .Z(n2198) );
  XOR2_X1 U3209 ( .A(n2651), .B(n2647), .Z(n2659) );
  XOR2_X1 U3058 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR2_X1 U3059 ( .A(n1953), .B(n1954), .Z(p6_S[38]) );
  XOR2_X1 U3130 ( .A(n2255), .B(n2254), .Z(n1951) );
  XOR2_X1 U3131 ( .A(n2253), .B(n2266), .Z(n2255) );
  XOR2_X1 U3132 ( .A(n2257), .B(n2258), .Z(n2266) );
  XOR2_X1 U2962 ( .A(n1489), .B(n1490), .Z(n1488) );
  XOR2_X1 U2965 ( .A(n1501), .B(n1502), .Z(n1500) );
  XOR2_X1 U3037 ( .A(n1805), .B(n1804), .Z(n1501) );
  XOR2_X1 U2851 ( .A(n906), .B(n905), .Z(n602) );
  XOR2_X1 U3056 ( .A(n1943), .B(n1944), .Z(n1942) );
  XOR2_X1 U3122 ( .A(n2201), .B(n2200), .Z(n1943) );
  XOR2_X1 U2933 ( .A(n1294), .B(n1293), .Z(n1298) );
  XOR2_X1 U3025 ( .A(n1761), .B(n1747), .Z(n1748) );
  MUX2_X1 U3033 ( .A(n1803), .B(n1804), .S(n1805), .Z(n1498) );
  XOR2_X1 U3100 ( .A(n2129), .B(n2131), .Z(n2161) );
  DFFR_X1 REGISTER4_q_reg_13_ ( .D(REGISTER4_n48), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[13]), .QN(n3773) );
  DFFR_X1 REG11_q_reg_9_ ( .D(REG11_n52), .CK(CLK), .RN(RST_n), .Q(reg2[9]), 
        .QN(n3691) );
  DFFR_X1 REG11_q_reg_6_ ( .D(REG11_n55), .CK(CLK), .RN(RST_n), .Q(reg2[6]), 
        .QN(n3687) );
  DFFR_X1 REG11_q_reg_4_ ( .D(REG11_n57), .CK(CLK), .RN(RST_n), .Q(reg2[4]), 
        .QN(n3685) );
  DFFR_X1 REG31_q_reg_9_ ( .D(REG31_n52), .CK(CLK), .RN(RST_n), .Q(reg4[9]), 
        .QN(n3681) );
  DFFR_X1 REG31_q_reg_6_ ( .D(REG31_n55), .CK(CLK), .RN(RST_n), .Q(reg4[6]), 
        .QN(n3678) );
  DFFR_X1 REG31_q_reg_0_ ( .D(REG31_n61), .CK(CLK), .RN(RST_n), .Q(reg4[0]), 
        .QN(n3670) );
  DFFR_X1 REGISTER2_q_reg_3_ ( .D(REGISTER2_n58), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[3]), .QN(n3718) );
  DFFR_X1 REG11_q_reg_7_ ( .D(REG11_n54), .CK(CLK), .RN(RST_n), .Q(reg2[7]), 
        .QN(n3688) );
  AOI22_X1 U1694 ( .A1(reg2[10]), .A2(n2326), .B1(n2324), .B2(n3693), .ZN(
        n2440) );
  AOI221_X1 U1693 ( .B1(n2328), .B2(reg2[11]), .C1(n2329), .C2(n3686), .A(
        n2440), .ZN(n2344) );
  AOI22_X1 U1692 ( .A1(reg2[13]), .A2(n2438), .B1(n2439), .B2(n3680), .ZN(
        n2431) );
  OAI221_X1 U1691 ( .B1(reg2[12]), .B2(n2429), .C1(n3690), .C2(n2430), .A(
        n2431), .ZN(n2432) );
  AOI22_X1 U1708 ( .A1(reg2[13]), .A2(n2456), .B1(n2457), .B2(n3680), .ZN(
        n2448) );
  AOI22_X1 U1699 ( .A1(reg2[12]), .A2(n2438), .B1(n2439), .B2(n3690), .ZN(
        n2449) );
  OAI221_X1 U1698 ( .B1(reg2[11]), .B2(n2429), .C1(n3686), .C2(n2430), .A(
        n2449), .ZN(n2436) );
  AOI22_X1 U1690 ( .A1(n2435), .A2(n2436), .B1(A1[13]), .B2(n2437), .ZN(n2346)
         );
  AOI222_X1 U1689 ( .A1(n2344), .A2(n2432), .B1(n2344), .B2(n2346), .C1(n2432), 
        .C2(n2346), .ZN(p11_C[53]) );
  AOI22_X1 U1688 ( .A1(reg2[11]), .A2(n2326), .B1(n2324), .B2(n3686), .ZN(
        n2433) );
  AOI221_X1 U1687 ( .B1(n2328), .B2(reg2[12]), .C1(n2329), .C2(n3690), .A(
        n2433), .ZN(n2342) );
  OAI221_X1 U1685 ( .B1(reg2[13]), .B2(n2429), .C1(n3680), .C2(n2430), .A(
        n2431), .ZN(n2341) );
  XNOR2_X1 U1661 ( .A(n2340), .B(n2341), .ZN(p11_S[54]) );
  XNOR2_X1 U1663 ( .A(n2343), .B(n2346), .ZN(n2345) );
  XNOR2_X1 U1662 ( .A(n2344), .B(n2345), .ZN(p11_S[53]) );
  AOI22_X1 U1710 ( .A1(reg2[10]), .A2(n2430), .B1(n2429), .B2(n3693), .ZN(
        n2458) );
  AOI221_X1 U1709 ( .B1(n2438), .B2(reg2[11]), .C1(n2439), .C2(n3686), .A(
        n2458), .ZN(n2452) );
  AOI22_X1 U1705 ( .A1(reg2[8]), .A2(n2326), .B1(n2324), .B2(n3683), .ZN(n2454) );
  AOI221_X1 U1704 ( .B1(n2328), .B2(reg2[9]), .C1(n2329), .C2(n3691), .A(n2454), .ZN(n2451) );
  OAI22_X1 U1701 ( .A1(n2450), .A2(n2451), .B1(n2452), .B2(n2349), .ZN(n2350)
         );
  AOI222_X1 U1695 ( .A1(n2442), .A2(n2443), .B1(n2442), .B2(n2348), .C1(n2443), 
        .C2(n2348), .ZN(p11_C[52]) );
  XNOR2_X1 U1754 ( .A(n2499), .B(n2500), .ZN(n2501) );
  AOI221_X1 U1752 ( .B1(n2456), .B2(reg2[10]), .C1(n2457), .C2(n3693), .A(
        n2516), .ZN(n2502) );
  OAI22_X1 U1739 ( .A1(n2499), .A2(n2500), .B1(n2501), .B2(n2502), .ZN(n2481)
         );
  AOI221_X1 U1735 ( .B1(n2456), .B2(reg2[11]), .C1(n2457), .C2(n3686), .A(
        n2496), .ZN(n2483) );
  AOI22_X1 U1734 ( .A1(reg2[8]), .A2(n2430), .B1(n2429), .B2(n3683), .ZN(n2495) );
  AOI221_X1 U1733 ( .B1(n2438), .B2(reg2[9]), .C1(n2439), .C2(n3691), .A(n2495), .ZN(n2494) );
  AOI22_X1 U1730 ( .A1(reg2[7]), .A2(n2328), .B1(n2329), .B2(n3688), .ZN(n2492) );
  OAI221_X1 U1729 ( .B1(reg2[6]), .B2(n2324), .C1(n3687), .C2(n2326), .A(n2492), .ZN(n2476) );
  XNOR2_X1 U1751 ( .A(n2501), .B(n2502), .ZN(n2488) );
  AOI22_X1 U1749 ( .A1(reg2[7]), .A2(n2430), .B1(n2429), .B2(n3688), .ZN(n2514) );
  AOI221_X1 U1748 ( .B1(n2438), .B2(reg2[8]), .C1(n2439), .C2(n3683), .A(n2514), .ZN(n2489) );
  XNOR2_X1 U1769 ( .A(n2521), .B(n2485), .ZN(n2522) );
  AOI22_X1 U1768 ( .A1(reg2[9]), .A2(n2456), .B1(n2457), .B2(n3691), .ZN(n2530) );
  OAI22_X1 U1758 ( .A1(n2521), .A2(n2485), .B1(n2522), .B2(n2523), .ZN(n2515)
         );
  XNOR2_X1 U1750 ( .A(n2515), .B(n2488), .ZN(n2490) );
  XNOR2_X1 U1747 ( .A(n2490), .B(n2489), .ZN(n2510) );
  AOI22_X1 U1746 ( .A1(reg2[5]), .A2(n2326), .B1(n2324), .B2(n3677), .ZN(n2512) );
  AOI22_X1 U1728 ( .A1(n2484), .A2(n2485), .B1(n2486), .B2(n2487), .ZN(n2359)
         );
  AOI222_X1 U1727 ( .A1(n2361), .A2(n2362), .B1(n2361), .B2(n2359), .C1(n2362), 
        .C2(n2359), .ZN(p11_C[49]) );
  AOI221_X1 U1721 ( .B1(n2456), .B2(reg2[12]), .C1(n2457), .C2(n3690), .A(
        n2474), .ZN(n2470) );
  AOI22_X1 U1718 ( .A1(reg2[9]), .A2(n2430), .B1(n2429), .B2(n3691), .ZN(n2469) );
  AOI221_X1 U1717 ( .B1(n2438), .B2(reg2[10]), .C1(n2439), .C2(n3693), .A(
        n2469), .ZN(n2463) );
  XNOR2_X1 U1716 ( .A(n2465), .B(n2463), .ZN(n2466) );
  AOI22_X1 U1715 ( .A1(reg2[8]), .A2(n2328), .B1(n2329), .B2(n3683), .ZN(n2468) );
  OAI221_X1 U1714 ( .B1(reg2[7]), .B2(n2324), .C1(n3688), .C2(n2326), .A(n2468), .ZN(n2460) );
  AOI22_X1 U1724 ( .A1(n2479), .A2(n2480), .B1(n2481), .B2(n2482), .ZN(n2357)
         );
  AOI22_X1 U1723 ( .A1(n2475), .A2(n2476), .B1(n2477), .B2(n2478), .ZN(n2358)
         );
  XNOR2_X1 U1666 ( .A(n2355), .B(n2356), .ZN(p11_S[50]) );
  XNOR2_X1 U1667 ( .A(n2359), .B(n2360), .ZN(p11_S[49]) );
  AOI22_X1 U1821 ( .A1(reg2[13]), .A2(n2601), .B1(n2602), .B2(n3680), .ZN(
        n2563) );
  NAND2_X1 U1775 ( .A1(n2534), .A2(n2537), .ZN(n2536) );
  AOI221_X1 U1792 ( .B1(n2456), .B2(reg2[8]), .C1(n2457), .C2(n3683), .A(n2564), .ZN(n2539) );
  AOI22_X1 U1786 ( .A1(reg2[6]), .A2(n2438), .B1(n2439), .B2(n3687), .ZN(n2556) );
  OAI221_X1 U1785 ( .B1(reg2[5]), .B2(n2429), .C1(n3677), .C2(n2430), .A(n2556), .ZN(n2542) );
  AOI22_X1 U1776 ( .A1(n2538), .A2(n2539), .B1(n2540), .B2(n2541), .ZN(n2507)
         );
  AOI22_X1 U1741 ( .A1(n2506), .A2(n2507), .B1(n2508), .B2(n2509), .ZN(n2366)
         );
  AOI22_X1 U1762 ( .A1(reg2[4]), .A2(n2326), .B1(n2324), .B2(n3685), .ZN(n2524) );
  AOI221_X1 U1761 ( .B1(n2328), .B2(reg2[5]), .C1(n2329), .C2(n3677), .A(n2524), .ZN(n2503) );
  AOI22_X1 U1765 ( .A1(reg2[6]), .A2(n2430), .B1(n2429), .B2(n3687), .ZN(n2527) );
  AOI221_X1 U1764 ( .B1(n2438), .B2(reg2[7]), .C1(n2439), .C2(n3688), .A(n2527), .ZN(n2504) );
  XNOR2_X1 U1763 ( .A(n2526), .B(n2504), .ZN(n2505) );
  AOI222_X1 U1740 ( .A1(n2365), .A2(n2366), .B1(n2365), .B2(n2363), .C1(n2366), 
        .C2(n2363), .ZN(p11_C[48]) );
  XNOR2_X1 U1760 ( .A(n2505), .B(n2503), .ZN(n2367) );
  XNOR2_X1 U1819 ( .A(n2600), .B(n2545), .ZN(n2555) );
  AOI22_X1 U1812 ( .A1(reg2[4]), .A2(n2430), .B1(n2429), .B2(n3685), .ZN(n2596) );
  AOI221_X1 U1811 ( .B1(n2438), .B2(reg2[5]), .C1(n2439), .C2(n3677), .A(n2596), .ZN(n2567) );
  AOI221_X1 U1817 ( .B1(n2456), .B2(reg2[7]), .C1(n2457), .C2(n3688), .A(n2599), .ZN(n2568) );
  XNOR2_X1 U1816 ( .A(n2555), .B(n2568), .ZN(n2597) );
  XNOR2_X1 U1813 ( .A(n2597), .B(n2554), .ZN(n2569) );
  AOI22_X1 U1780 ( .A1(n2547), .A2(n2548), .B1(n2549), .B2(n2550), .ZN(n2369)
         );
  AOI22_X1 U1795 ( .A1(reg2[4]), .A2(n2328), .B1(n2329), .B2(n3685), .ZN(n2566) );
  OAI221_X1 U1794 ( .B1(reg2[3]), .B2(n2324), .C1(n3669), .C2(n2326), .A(n2566), .ZN(n2544) );
  AOI22_X1 U1779 ( .A1(n2543), .A2(n2544), .B1(n2545), .B2(n2546), .ZN(n2370)
         );
  XNOR2_X1 U1669 ( .A(n2367), .B(n2368), .ZN(p11_S[47]) );
  XNOR2_X1 U1810 ( .A(n2569), .B(n2567), .ZN(n2575) );
  AOI22_X1 U1835 ( .A1(reg2[13]), .A2(n2334), .B1(A1[1]), .B2(n3680), .ZN(
        n2625) );
  AOI22_X1 U1833 ( .A1(reg2[12]), .A2(n2601), .B1(n2602), .B2(n3690), .ZN(
        n2624) );
  AOI22_X1 U1829 ( .A1(reg2[6]), .A2(n2456), .B1(n2457), .B2(n3687), .ZN(n2620) );
  AOI22_X1 U1843 ( .A1(reg2[3]), .A2(n2430), .B1(n2429), .B2(n3669), .ZN(n2629) );
  AOI221_X1 U1842 ( .B1(n2438), .B2(reg2[4]), .C1(n2439), .C2(n3685), .A(n2629), .ZN(n2573) );
  AOI22_X1 U1841 ( .A1(reg2[1]), .A2(n2326), .B1(n2324), .B2(n3684), .ZN(n2628) );
  NOR2_X1 U1809 ( .A1(n2573), .A2(n2574), .ZN(n2591) );
  XNOR2_X1 U1808 ( .A(n2577), .B(n2591), .ZN(n2586) );
  XNOR2_X1 U1805 ( .A(n2586), .B(n2576), .ZN(n2570) );
  AOI22_X1 U1804 ( .A1(reg2[3]), .A2(n2328), .B1(n2329), .B2(n3669), .ZN(n2585) );
  OAI221_X1 U1803 ( .B1(reg2[2]), .B2(n2324), .C1(n3692), .C2(n2326), .A(n2585), .ZN(n2571) );
  OAI21_X1 U1797 ( .B1(n2573), .B2(n2574), .A(n2570), .ZN(n2572) );
  OAI21_X1 U1796 ( .B1(n2570), .B2(n2571), .A(n2572), .ZN(n2374) );
  AOI222_X1 U1783 ( .A1(n2373), .A2(n2374), .B1(n2373), .B2(n2371), .C1(n2374), 
        .C2(n2371), .ZN(p11_C[46]) );
  AOI221_X1 U1851 ( .B1(n2456), .B2(reg2[5]), .C1(n2457), .C2(n3677), .A(n2637), .ZN(n2613) );
  AOI221_X1 U1862 ( .B1(n2601), .B2(reg2[11]), .C1(n2602), .C2(n3686), .A(
        n2643), .ZN(n2641) );
  NAND2_X1 U2038 ( .A1(A1[0]), .A2(A1[1]), .ZN(n2337) );
  AOI22_X1 U1861 ( .A1(reg2[13]), .A2(n2334), .B1(n2335), .B2(n3680), .ZN(
        n2642) );
  OAI21_X1 U1860 ( .B1(reg2[12]), .B2(n2332), .A(n2642), .ZN(n2615) );
  XNOR2_X1 U1859 ( .A(n2641), .B(n2615), .ZN(n2616) );
  AOI221_X1 U1857 ( .B1(n2531), .B2(reg2[9]), .C1(n2532), .C2(n3691), .A(n2640), .ZN(n2618) );
  XNOR2_X1 U1853 ( .A(n2638), .B(n2612), .ZN(n2614) );
  XNOR2_X1 U1839 ( .A(n2573), .B(n2574), .ZN(n2619) );
  OAI21_X1 U1826 ( .B1(n2615), .B2(n2616), .A(n2617), .ZN(n2582) );
  XNOR2_X1 U1671 ( .A(n2377), .B(n2378), .ZN(n2375) );
  AOI22_X1 U1799 ( .A1(n2578), .A2(n2579), .B1(n2580), .B2(n2581), .ZN(n2376)
         );
  AOI221_X1 U1876 ( .B1(n2456), .B2(reg2[4]), .C1(n2457), .C2(n3685), .A(n2663), .ZN(n2645) );
  OAI22_X1 U1886 ( .A1(reg2[11]), .A2(n2332), .B1(reg2[12]), .B2(n2337), .ZN(
        n2668) );
  AOI21_X1 U1885 ( .B1(reg2[12]), .B2(n2334), .A(n2668), .ZN(n2634) );
  AOI22_X1 U1847 ( .A1(reg2[0]), .A2(n2326), .B1(n2324), .B2(n3689), .ZN(n2630) );
  AOI22_X1 U1849 ( .A1(reg2[2]), .A2(n2430), .B1(n2429), .B2(n3692), .ZN(n2632) );
  AOI221_X1 U1848 ( .B1(n2438), .B2(reg2[3]), .C1(n2439), .C2(n3669), .A(n2632), .ZN(n2605) );
  AOI222_X1 U1824 ( .A1(n2381), .A2(n2382), .B1(n2381), .B2(n2379), .C1(n2382), 
        .C2(n2379), .ZN(p11_C[44]) );
  AOI221_X1 U1913 ( .B1(n2601), .B2(reg2[9]), .C1(n2602), .C2(n3691), .A(n2694), .ZN(n2670) );
  OAI22_X1 U1912 ( .A1(reg2[11]), .A2(n2337), .B1(reg2[10]), .B2(n2332), .ZN(
        n2693) );
  AOI21_X1 U1911 ( .B1(reg2[11]), .B2(n2334), .A(n2693), .ZN(n2671) );
  AOI22_X1 U1891 ( .A1(reg2[1]), .A2(n2430), .B1(n2429), .B2(n3684), .ZN(n2673) );
  AOI221_X1 U1890 ( .B1(n2438), .B2(reg2[2]), .C1(n2439), .C2(n3692), .A(n2673), .ZN(n2649) );
  XNOR2_X1 U1845 ( .A(n2606), .B(n2604), .ZN(n2383) );
  XNOR2_X1 U1910 ( .A(n2670), .B(n2671), .ZN(n2691) );
  AOI221_X1 U1927 ( .B1(n2531), .B2(reg2[6]), .C1(n2532), .C2(n3687), .A(n2700), .ZN(n2686) );
  AOI221_X1 U1896 ( .B1(n2456), .B2(reg2[3]), .C1(n2457), .C2(n3669), .A(n2682), .ZN(n2652) );
  AOI22_X1 U1894 ( .A1(reg2[0]), .A2(n2430), .B1(n2429), .B2(n3689), .ZN(n2680) );
  AOI221_X1 U1893 ( .B1(n2438), .B2(reg2[1]), .C1(n2439), .C2(n3684), .A(n2680), .ZN(n2653) );
  XNOR2_X1 U1898 ( .A(n2657), .B(n2656), .ZN(n2681) );
  XNOR2_X1 U1895 ( .A(n2681), .B(n2652), .ZN(n2654) );
  AOI221_X1 U1932 ( .B1(n2456), .B2(reg2[2]), .C1(n2457), .C2(n3692), .A(n2704), .ZN(n2678) );
  AOI22_X1 U1939 ( .A1(reg2[9]), .A2(n2334), .B1(n2335), .B2(n3691), .ZN(n2720) );
  OAI21_X1 U1938 ( .B1(reg2[8]), .B2(n2332), .A(n2720), .ZN(n2702) );
  AOI221_X1 U1918 ( .B1(n2438), .B2(reg2[0]), .C1(n2439), .C2(n3689), .A(n2697), .ZN(n2675) );
  AOI222_X1 U1892 ( .A1(n2393), .A2(n2394), .B1(n2393), .B2(n2391), .C1(n2394), 
        .C2(n2391), .ZN(p11_C[41]) );
  AOI22_X1 U1966 ( .A1(reg2[8]), .A2(n2334), .B1(n2335), .B2(n3683), .ZN(n2736) );
  OAI21_X1 U1965 ( .B1(reg2[7]), .B2(n2332), .A(n2736), .ZN(n2722) );
  NAND2_X1 U1942 ( .A1(n2722), .A2(n2723), .ZN(n2719) );
  AOI221_X1 U1935 ( .B1(n2456), .B2(reg2[1]), .C1(n2457), .C2(n3684), .A(n2717), .ZN(n2706) );
  XNOR2_X1 U1964 ( .A(n2723), .B(n2722), .ZN(n2715) );
  XNOR2_X1 U1963 ( .A(n2735), .B(n2715), .ZN(n2716) );
  AOI221_X1 U1986 ( .B1(n2601), .B2(reg2[5]), .C1(n2602), .C2(n3677), .A(n2751), .ZN(n2727) );
  OAI22_X1 U1985 ( .A1(reg2[6]), .A2(n2332), .B1(reg2[7]), .B2(n2337), .ZN(
        n2750) );
  AOI21_X1 U1984 ( .B1(n2334), .B2(reg2[7]), .A(n2750), .ZN(n2728) );
  AOI221_X1 U1981 ( .B1(n2531), .B2(reg2[3]), .C1(n2532), .C2(n3669), .A(n2749), .ZN(n2729) );
  AOI222_X1 U1949 ( .A1(n2727), .A2(n2728), .B1(n2727), .B2(n2729), .C1(n2728), 
        .C2(n2729), .ZN(n2726) );
  AOI22_X1 U2010 ( .A1(reg2[5]), .A2(n2334), .B1(n2335), .B2(n3677), .ZN(n2761) );
  OAI21_X1 U2009 ( .B1(reg2[4]), .B2(n2332), .A(n2761), .ZN(n2413) );
  AOI22_X1 U1977 ( .A1(n3677), .A2(n2746), .B1(n3669), .B2(n2747), .ZN(n2745)
         );
  OAI221_X1 U1976 ( .B1(n2339), .B2(n3687), .C1(n2337), .C2(reg2[6]), .A(n2745), .ZN(n2744) );
  AOI221_X1 U1975 ( .B1(n3685), .B2(n2602), .C1(reg2[4]), .C2(n2601), .A(n2744), .ZN(n2740) );
  AOI221_X1 U1973 ( .B1(n2740), .B2(n3669), .C1(n2740), .C2(n2562), .A(n2741), 
        .ZN(n2405) );
  XNOR2_X1 U1983 ( .A(n2727), .B(n2728), .ZN(n2748) );
  XNOR2_X1 U1980 ( .A(n2748), .B(n2729), .ZN(n2408) );
  AOI22_X1 U2018 ( .A1(reg2[4]), .A2(n2334), .B1(n2335), .B2(n3685), .ZN(n2764) );
  OAI21_X1 U2017 ( .B1(reg2[3]), .B2(n2332), .A(n2764), .ZN(n2420) );
  NAND2_X1 U1682 ( .A1(n2419), .A2(n2420), .ZN(n2418) );
  XNOR2_X1 U1681 ( .A(n2417), .B(n2418), .ZN(n2416) );
  XNOR2_X1 U2014 ( .A(n2420), .B(n2419), .ZN(n2422) );
  AOI221_X1 U2032 ( .B1(n2602), .B2(n3684), .C1(n2601), .C2(reg2[1]), .A(n2769), .ZN(n2425) );
  AOI22_X1 U2030 ( .A1(reg2[3]), .A2(n2334), .B1(n2335), .B2(n3669), .ZN(n2768) );
  OAI21_X1 U2029 ( .B1(reg2[2]), .B2(n2332), .A(n2768), .ZN(n2767) );
  AOI22_X1 U1659 ( .A1(reg2[1]), .A2(n2334), .B1(n2335), .B2(n3684), .ZN(n2333) );
  OAI21_X1 U1658 ( .B1(reg2[0]), .B2(n2332), .A(n2333), .ZN(
        p11_final_product1[1]) );
  OAI221_X1 U1660 ( .B1(reg2[0]), .B2(n2337), .C1(n3689), .C2(n2339), .A(n2332), .ZN(p11_final_product1[0]) );
  NOR2_X1 U2027 ( .A1(n2425), .A2(n2426), .ZN(p11_C[33]) );
  OAI211_X1 U2006 ( .C1(n2417), .C2(n2415), .A(n2420), .B(n2419), .ZN(n2758)
         );
  NAND2_X1 U2005 ( .A1(n2417), .A2(n2415), .ZN(n2759) );
  NAND2_X1 U2004 ( .A1(n2758), .A2(n2759), .ZN(p11_C[35]) );
  NAND2_X1 U1680 ( .A1(n2413), .A2(n2414), .ZN(n2412) );
  XNOR2_X1 U1678 ( .A(n2409), .B(n2410), .ZN(p11_S[36]) );
  AOI222_X1 U1971 ( .A1(n2407), .A2(n2408), .B1(n2407), .B2(n2739), .C1(n2408), 
        .C2(n2739), .ZN(p11_C[37]) );
  AOI222_X1 U1844 ( .A1(n2385), .A2(n2386), .B1(n2385), .B2(n2383), .C1(n2386), 
        .C2(n2383), .ZN(p11_C[43]) );
  XNOR2_X1 U1670 ( .A(n2371), .B(n2372), .ZN(p11_S[46]) );
  AOI222_X1 U1798 ( .A1(n2377), .A2(n2378), .B1(n2377), .B2(n2376), .C1(n2378), 
        .C2(n2376), .ZN(p11_C[45]) );
  XNOR2_X1 U1668 ( .A(n2363), .B(n2364), .ZN(p11_S[48]) );
  AOI222_X1 U1759 ( .A1(n2369), .A2(n2370), .B1(n2369), .B2(n2367), .C1(n2370), 
        .C2(n2367), .ZN(p11_C[47]) );
  AOI222_X1 U1713 ( .A1(n2357), .A2(n2358), .B1(n2357), .B2(n2355), .C1(n2358), 
        .C2(n2355), .ZN(p11_C[50]) );
  XNOR2_X1 U1703 ( .A(n2450), .B(n2451), .ZN(n2351) );
  XNOR2_X1 U1665 ( .A(n2351), .B(n2352), .ZN(p11_S[51]) );
  XNOR2_X1 U1664 ( .A(n2347), .B(n2348), .ZN(p11_S[52]) );
  AOI222_X1 U1702 ( .A1(n2353), .A2(n2354), .B1(n2353), .B2(n2351), .C1(n2354), 
        .C2(n2351), .ZN(p11_C[51]) );
  AOI22_X1 U1656 ( .A1(reg2[13]), .A2(n2328), .B1(n2329), .B2(n3680), .ZN(
        n2327) );
  OAI221_X1 U1655 ( .B1(reg2[12]), .B2(n2324), .C1(n3690), .C2(n2326), .A(
        n2327), .ZN(p11_final_product2_26_) );
  NOR2_X1 U60 ( .A1(n2331), .A2(n2328), .ZN(n523) );
  NOR2_X1 U1077 ( .A1(n3694), .A2(n3725), .ZN(n1431) );
  OAI21_X1 U1075 ( .B1(reg2_reg[11]), .B2(reg2_reg[12]), .A(n1426), .ZN(n1758)
         );
  AOI22_X1 U890 ( .A1(B1[11]), .A2(n1426), .B1(n1424), .B2(n1534), .ZN(n1533)
         );
  AOI221_X1 U889 ( .B1(n1428), .B2(B1[12]), .C1(n1429), .C2(n1425), .A(n1533), 
        .ZN(n1442) );
  OAI21_X1 U1126 ( .B1(reg2_reg[9]), .B2(reg2_reg[10]), .A(n1530), .ZN(n1796)
         );
  AOI22_X1 U894 ( .A1(B1[13]), .A2(n1538), .B1(n1539), .B2(n1430), .ZN(n1531)
         );
  OAI221_X1 U893 ( .B1(B1[12]), .B2(n1529), .C1(n1425), .C2(n1530), .A(n1531), 
        .ZN(n1532) );
  OAI221_X1 U887 ( .B1(B1[13]), .B2(n1529), .C1(n1430), .C2(n1530), .A(n1531), 
        .ZN(n1441) );
  AOI22_X1 U860 ( .A1(B1[13]), .A2(n1428), .B1(n1429), .B2(n1430), .ZN(n1427)
         );
  OAI221_X1 U859 ( .B1(B1[12]), .B2(n1424), .C1(n1425), .C2(n1426), .A(n1427), 
        .ZN(p7_final_product2_26_) );
  AOI22_X1 U896 ( .A1(B1[10]), .A2(n1426), .B1(n1424), .B2(n1541), .ZN(n1540)
         );
  AOI221_X1 U895 ( .B1(n1428), .B2(B1[11]), .C1(n1429), .C2(n1534), .A(n1540), 
        .ZN(n1444) );
  OAI21_X1 U1162 ( .B1(reg2_reg[7]), .B2(reg2_reg[8]), .A(n1547), .ZN(n1831)
         );
  AOI22_X1 U910 ( .A1(B1[13]), .A2(n1556), .B1(n1557), .B2(n1430), .ZN(n1548)
         );
  OAI221_X1 U899 ( .B1(B1[13]), .B2(n1546), .C1(n1430), .C2(n1547), .A(n1548), 
        .ZN(n1545) );
  AOI22_X1 U901 ( .A1(B1[12]), .A2(n1538), .B1(n1539), .B2(n1425), .ZN(n1549)
         );
  OAI221_X1 U900 ( .B1(B1[11]), .B2(n1529), .C1(n1534), .C2(n1530), .A(n1549), 
        .ZN(n1536) );
  AOI22_X1 U892 ( .A1(n1535), .A2(n1536), .B1(reg2_reg[13]), .B2(n1537), .ZN(
        n1446) );
  XNOR2_X1 U866 ( .A(n1443), .B(n1446), .ZN(n1445) );
  XNOR2_X1 U865 ( .A(n1444), .B(n1445), .ZN(p7_S[53]) );
  OAI221_X1 U909 ( .B1(B1[12]), .B2(n1546), .C1(n1425), .C2(n1547), .A(n1548), 
        .ZN(n1449) );
  AOI22_X1 U912 ( .A1(B1[10]), .A2(n1530), .B1(n1529), .B2(n1541), .ZN(n1558)
         );
  AOI221_X1 U911 ( .B1(n1538), .B2(B1[11]), .C1(n1539), .C2(n1534), .A(n1558), 
        .ZN(n1552) );
  AOI221_X1 U906 ( .B1(n1428), .B2(B1[9]), .C1(n1429), .C2(n1553), .A(n1554), 
        .ZN(n1551) );
  OAI22_X1 U903 ( .A1(n1550), .A2(n1551), .B1(n1552), .B2(n1449), .ZN(n1450)
         );
  AOI222_X1 U897 ( .A1(n1542), .A2(n1543), .B1(n1542), .B2(n1448), .C1(n1543), 
        .C2(n1448), .ZN(p7_C[52]) );
  XNOR2_X1 U905 ( .A(n1550), .B(n1551), .ZN(n1451) );
  AOI22_X1 U920 ( .A1(B1[9]), .A2(n1530), .B1(n1529), .B2(n1553), .ZN(n1569)
         );
  AOI221_X1 U919 ( .B1(n1538), .B2(B1[10]), .C1(n1539), .C2(n1541), .A(n1569), 
        .ZN(n1563) );
  OAI21_X1 U1203 ( .B1(reg2_reg[6]), .B2(reg2_reg[5]), .A(n1572), .ZN(n1854)
         );
  AOI22_X1 U940 ( .A1(B1[13]), .A2(n1597), .B1(n1598), .B2(n1430), .ZN(n1573)
         );
  OAI221_X1 U922 ( .B1(B1[13]), .B2(n1571), .C1(n1430), .C2(n1572), .A(n1573), 
        .ZN(n1564) );
  AOI22_X1 U924 ( .A1(B1[11]), .A2(n1547), .B1(n1546), .B2(n1534), .ZN(n1574)
         );
  AOI221_X1 U923 ( .B1(n1556), .B2(B1[12]), .C1(n1557), .C2(n1425), .A(n1574), 
        .ZN(n1570) );
  XNOR2_X1 U921 ( .A(n1570), .B(n1564), .ZN(n1565) );
  XNOR2_X1 U918 ( .A(n1565), .B(n1563), .ZN(n1566) );
  OAI221_X1 U916 ( .B1(B1[7]), .B2(n1424), .C1(n1567), .C2(n1426), .A(n1568), 
        .ZN(n1560) );
  OAI221_X1 U939 ( .B1(B1[12]), .B2(n1571), .C1(n1425), .C2(n1572), .A(n1573), 
        .ZN(n1561) );
  AOI22_X1 U913 ( .A1(n1559), .A2(n1560), .B1(n1561), .B2(n1562), .ZN(n1454)
         );
  XNOR2_X1 U868 ( .A(n1451), .B(n1452), .ZN(p7_S[51]) );
  AOI22_X1 U959 ( .A1(B1[11]), .A2(n1572), .B1(n1571), .B2(n1534), .ZN(n1620)
         );
  AOI221_X1 U958 ( .B1(n1597), .B2(B1[12]), .C1(n1598), .C2(n1425), .A(n1620), 
        .ZN(n1599) );
  OAI21_X1 U1228 ( .B1(reg2_reg[3]), .B2(reg2_reg[4]), .A(n1618), .ZN(n1863)
         );
  AOI22_X1 U973 ( .A1(B1[13]), .A2(n1631), .B1(n1632), .B2(n1430), .ZN(n1619)
         );
  OAI221_X1 U957 ( .B1(B1[13]), .B2(n1617), .C1(n1430), .C2(n1618), .A(n1619), 
        .ZN(n1600) );
  XNOR2_X1 U956 ( .A(n1599), .B(n1600), .ZN(n1601) );
  AOI22_X1 U955 ( .A1(B1[9]), .A2(n1547), .B1(n1546), .B2(n1553), .ZN(n1616)
         );
  AOI221_X1 U954 ( .B1(n1556), .B2(B1[10]), .C1(n1557), .C2(n1541), .A(n1616), 
        .ZN(n1602) );
  OAI22_X1 U941 ( .A1(n1599), .A2(n1600), .B1(n1601), .B2(n1602), .ZN(n1581)
         );
  AOI22_X1 U938 ( .A1(B1[10]), .A2(n1547), .B1(n1546), .B2(n1541), .ZN(n1596)
         );
  AOI221_X1 U937 ( .B1(n1556), .B2(B1[11]), .C1(n1557), .C2(n1534), .A(n1596), 
        .ZN(n1583) );
  AOI22_X1 U926 ( .A1(n1579), .A2(n1580), .B1(n1581), .B2(n1582), .ZN(n1457)
         );
  AOI221_X1 U935 ( .B1(n1538), .B2(B1[9]), .C1(n1539), .C2(n1553), .A(n1595), 
        .ZN(n1594) );
  AOI22_X1 U932 ( .A1(B1[7]), .A2(n1428), .B1(n1429), .B2(n1567), .ZN(n1592)
         );
  OAI221_X1 U931 ( .B1(B1[6]), .B2(n1424), .C1(n1591), .C2(n1426), .A(n1592), 
        .ZN(n1576) );
  AOI22_X1 U925 ( .A1(n1575), .A2(n1576), .B1(n1577), .B2(n1578), .ZN(n1458)
         );
  AOI222_X1 U915 ( .A1(n1457), .A2(n1458), .B1(n1457), .B2(n1455), .C1(n1458), 
        .C2(n1455), .ZN(p7_C[50]) );
  AOI22_X1 U975 ( .A1(B1[10]), .A2(n1572), .B1(n1571), .B2(n1541), .ZN(n1633)
         );
  AOI221_X1 U974 ( .B1(n1597), .B2(B1[11]), .C1(n1598), .C2(n1534), .A(n1633), 
        .ZN(n1621) );
  OAI221_X1 U972 ( .B1(B1[12]), .B2(n1617), .C1(n1425), .C2(n1618), .A(n1619), 
        .ZN(n1585) );
  XNOR2_X1 U971 ( .A(n1621), .B(n1585), .ZN(n1622) );
  AOI22_X1 U970 ( .A1(B1[9]), .A2(n1556), .B1(n1557), .B2(n1553), .ZN(n1630)
         );
  OAI22_X1 U960 ( .A1(n1621), .A2(n1585), .B1(n1622), .B2(n1623), .ZN(n1615)
         );
  XNOR2_X1 U953 ( .A(n1601), .B(n1602), .ZN(n1588) );
  XNOR2_X1 U952 ( .A(n1615), .B(n1588), .ZN(n1590) );
  AOI22_X1 U951 ( .A1(B1[7]), .A2(n1530), .B1(n1529), .B2(n1567), .ZN(n1614)
         );
  XNOR2_X1 U949 ( .A(n1590), .B(n1589), .ZN(n1610) );
  AOI22_X1 U930 ( .A1(n1584), .A2(n1585), .B1(n1586), .B2(n1587), .ZN(n1459)
         );
  XNOR2_X1 U870 ( .A(n1459), .B(n1460), .ZN(p7_S[49]) );
  OAI21_X1 U1254 ( .B1(reg2_reg[1]), .B2(reg2_reg[2]), .A(n1662), .ZN(n1872)
         );
  AOI22_X1 U1023 ( .A1(B1[13]), .A2(n1698), .B1(n1699), .B2(n1430), .ZN(n1663)
         );
  OAI221_X1 U993 ( .B1(B1[13]), .B2(n1661), .C1(n1430), .C2(n1662), .A(n1663), 
        .ZN(n1637) );
  AOI22_X1 U992 ( .A1(B1[12]), .A2(n1631), .B1(n1632), .B2(n1425), .ZN(n1660)
         );
  OAI221_X1 U991 ( .B1(B1[11]), .B2(n1617), .C1(n1534), .C2(n1618), .A(n1660), 
        .ZN(n1659) );
  AOI22_X1 U990 ( .A1(B1[10]), .A2(n1597), .B1(n1598), .B2(n1541), .ZN(n1658)
         );
  OAI221_X1 U989 ( .B1(B1[9]), .B2(n1571), .C1(n1553), .C2(n1572), .A(n1658), 
        .ZN(n1635) );
  NAND2_X1 U977 ( .A1(n1634), .A2(n1637), .ZN(n1636) );
  OAI21_X1 U976 ( .B1(n1634), .B2(n1635), .A(n1636), .ZN(n1628) );
  AOI22_X1 U995 ( .A1(B1[7]), .A2(n1547), .B1(n1546), .B2(n1567), .ZN(n1664)
         );
  AOI22_X1 U988 ( .A1(B1[6]), .A2(n1538), .B1(n1539), .B2(n1591), .ZN(n1656)
         );
  AOI22_X1 U978 ( .A1(n1638), .A2(n1639), .B1(n1640), .B2(n1641), .ZN(n1607)
         );
  AOI22_X1 U943 ( .A1(n1606), .A2(n1607), .B1(n1608), .B2(n1609), .ZN(n1466)
         );
  AOI22_X1 U964 ( .A1(B1[4]), .A2(n1426), .B1(n1424), .B2(n1625), .ZN(n1624)
         );
  AOI22_X1 U967 ( .A1(B1[6]), .A2(n1530), .B1(n1529), .B2(n1591), .ZN(n1627)
         );
  AOI221_X1 U966 ( .B1(n1538), .B2(B1[7]), .C1(n1539), .C2(n1567), .A(n1627), 
        .ZN(n1604) );
  XNOR2_X1 U965 ( .A(n1626), .B(n1604), .ZN(n1605) );
  XNOR2_X1 U962 ( .A(n1605), .B(n1603), .ZN(n1467) );
  AOI221_X1 U1016 ( .B1(n1597), .B2(B1[9]), .C1(n1598), .C2(n1553), .A(n1695), 
        .ZN(n1654) );
  OAI221_X1 U1022 ( .B1(B1[12]), .B2(n1661), .C1(n1425), .C2(n1662), .A(n1663), 
        .ZN(n1645) );
  AOI221_X1 U1024 ( .B1(n1631), .B2(B1[11]), .C1(n1632), .C2(n1534), .A(n1700), 
        .ZN(n1697) );
  XNOR2_X1 U1021 ( .A(n1697), .B(n1645), .ZN(n1655) );
  AOI22_X1 U1014 ( .A1(B1[4]), .A2(n1530), .B1(n1529), .B2(n1625), .ZN(n1693)
         );
  AOI22_X1 U1020 ( .A1(B1[6]), .A2(n1547), .B1(n1546), .B2(n1591), .ZN(n1696)
         );
  XNOR2_X1 U1018 ( .A(n1655), .B(n1668), .ZN(n1694) );
  XNOR2_X1 U1015 ( .A(n1694), .B(n1654), .ZN(n1669) );
  AOI22_X1 U982 ( .A1(n1647), .A2(n1648), .B1(n1649), .B2(n1650), .ZN(n1469)
         );
  AOI22_X1 U997 ( .A1(B1[4]), .A2(n1428), .B1(n1429), .B2(n1625), .ZN(n1666)
         );
  OAI221_X1 U996 ( .B1(B1[3]), .B2(n1424), .C1(n1665), .C2(n1426), .A(n1666), 
        .ZN(n1644) );
  AOI22_X1 U981 ( .A1(n1643), .A2(n1644), .B1(n1645), .B2(n1646), .ZN(n1470)
         );
  XNOR2_X1 U872 ( .A(n1467), .B(n1468), .ZN(p7_S[47]) );
  XNOR2_X1 U1012 ( .A(n1669), .B(n1667), .ZN(n1675) );
  AOI22_X1 U1039 ( .A1(B1[7]), .A2(n1572), .B1(n1571), .B2(n1567), .ZN(n1721)
         );
  NAND2_X1 U1246 ( .A1(n3716), .A2(reg2_reg[0]), .ZN(n1439) );
  AOI22_X1 U1037 ( .A1(B1[13]), .A2(n1434), .B1(reg2_reg[1]), .B2(n1430), .ZN(
        n1701) );
  AOI22_X1 U1035 ( .A1(B1[11]), .A2(n1662), .B1(n1661), .B2(n1534), .ZN(n1720)
         );
  AOI221_X1 U1034 ( .B1(n1698), .B2(B1[12]), .C1(n1699), .C2(n1425), .A(n1720), 
        .ZN(n1719) );
  OAI221_X1 U1032 ( .B1(B1[9]), .B2(n1617), .C1(n1553), .C2(n1618), .A(n1718), 
        .ZN(n1704) );
  AOI22_X1 U1031 ( .A1(B1[6]), .A2(n1556), .B1(n1557), .B2(n1591), .ZN(n1716)
         );
  AOI22_X1 U1007 ( .A1(n1686), .A2(n1687), .B1(n1688), .B2(n1689), .ZN(n1676)
         );
  OAI22_X1 U1026 ( .A1(n1701), .A2(n1702), .B1(n1703), .B2(n1704), .ZN(n1692)
         );
  AOI22_X1 U1044 ( .A1(B1[3]), .A2(n1530), .B1(n1529), .B2(n1665), .ZN(n1723)
         );
  AOI22_X1 U1042 ( .A1(B1[1]), .A2(n1426), .B1(n1424), .B2(n1436), .ZN(n1722)
         );
  NOR2_X1 U1011 ( .A1(n1673), .A2(n1674), .ZN(n1691) );
  XNOR2_X1 U1010 ( .A(n1677), .B(n1691), .ZN(n1685) );
  XNOR2_X1 U1006 ( .A(n1685), .B(n1676), .ZN(n1670) );
  AOI22_X1 U1005 ( .A1(B1[3]), .A2(n1428), .B1(n1429), .B2(n1665), .ZN(n1684)
         );
  OAI21_X1 U999 ( .B1(n1673), .B2(n1674), .A(n1670), .ZN(n1672) );
  OAI21_X1 U998 ( .B1(n1670), .B2(n1671), .A(n1672), .ZN(n1474) );
  AOI222_X1 U985 ( .A1(n1473), .A2(n1474), .B1(n1473), .B2(n1471), .C1(n1474), 
        .C2(n1471), .ZN(p7_C[46]) );
  AOI22_X1 U1062 ( .A1(B1[7]), .A2(n1597), .B1(n1598), .B2(n1567), .ZN(n1739)
         );
  OAI221_X1 U1061 ( .B1(B1[6]), .B2(n1571), .C1(n1591), .C2(n1572), .A(n1739), 
        .ZN(n1712) );
  OAI221_X1 U1050 ( .B1(B1[4]), .B2(n1546), .C1(n1625), .C2(n1547), .A(n1733), 
        .ZN(n1713) );
  AOI221_X1 U1058 ( .B1(n1698), .B2(B1[11]), .C1(n1699), .C2(n1534), .A(n1738), 
        .ZN(n1736) );
  NAND2_X1 U1247 ( .A1(reg2_reg[1]), .A2(n3723), .ZN(n1432) );
  NAND2_X1 U1244 ( .A1(reg2_reg[0]), .A2(reg2_reg[1]), .ZN(n1437) );
  AOI22_X1 U1056 ( .A1(B1[13]), .A2(n1434), .B1(n1435), .B2(n1430), .ZN(n1737)
         );
  OAI21_X1 U1055 ( .B1(B1[12]), .B2(n1432), .A(n1737), .ZN(n1724) );
  XNOR2_X1 U1054 ( .A(n1736), .B(n1724), .ZN(n1726) );
  AOI22_X1 U1053 ( .A1(B1[9]), .A2(n1631), .B1(n1632), .B2(n1553), .ZN(n1735)
         );
  XNOR2_X1 U1040 ( .A(n1673), .B(n1674), .ZN(n1715) );
  XNOR2_X1 U1029 ( .A(n1711), .B(n1682), .ZN(n1481) );
  XNOR2_X1 U874 ( .A(n1477), .B(n1478), .ZN(n1475) );
  XNOR2_X1 U1049 ( .A(n1714), .B(n1713), .ZN(n1708) );
  AOI221_X1 U1084 ( .B1(n1597), .B2(B1[6]), .C1(n1598), .C2(n1591), .A(n1765), 
        .ZN(n1741) );
  AOI22_X1 U1079 ( .A1(B1[3]), .A2(n1547), .B1(n1546), .B2(n1665), .ZN(n1762)
         );
  OAI22_X1 U1090 ( .A1(B1[11]), .A2(n1432), .B1(B1[12]), .B2(n1437), .ZN(n1768) );
  AOI21_X1 U1089 ( .B1(B1[12]), .B2(n1434), .A(n1768), .ZN(n1730) );
  AOI22_X1 U1082 ( .A1(B1[7]), .A2(n1618), .B1(n1617), .B2(n1567), .ZN(n1764)
         );
  XNOR2_X1 U1080 ( .A(n1763), .B(n1731), .ZN(n1743) );
  AOI22_X1 U1048 ( .A1(B1[0]), .A2(n1426), .B1(n1424), .B2(n1438), .ZN(n1727)
         );
  XNOR2_X1 U1063 ( .A(n1709), .B(n1706), .ZN(n1728) );
  XNOR2_X1 U1046 ( .A(n1707), .B(n1705), .ZN(n1483) );
  AOI22_X1 U1093 ( .A1(B1[1]), .A2(n1530), .B1(n1529), .B2(n1436), .ZN(n1772)
         );
  AOI221_X1 U1116 ( .B1(n1698), .B2(B1[9]), .C1(n1699), .C2(n1553), .A(n1792), 
        .ZN(n1769) );
  OAI22_X1 U1115 ( .A1(B1[11]), .A2(n1437), .B1(B1[10]), .B2(n1432), .ZN(n1791) );
  AOI21_X1 U1114 ( .B1(B1[11]), .B2(n1434), .A(n1791), .ZN(n1770) );
  AOI22_X1 U1112 ( .A1(B1[6]), .A2(n1618), .B1(n1617), .B2(n1591), .ZN(n1790)
         );
  XNOR2_X1 U876 ( .A(n1483), .B(n1484), .ZN(p7_S[43]) );
  XNOR2_X1 U1110 ( .A(n1789), .B(n1771), .ZN(n1752) );
  AOI22_X1 U1102 ( .A1(B1[4]), .A2(n1572), .B1(n1571), .B2(n1625), .ZN(n1781)
         );
  AOI22_X1 U1132 ( .A1(B1[3]), .A2(n1572), .B1(n1571), .B2(n1665), .ZN(n1799)
         );
  NOR2_X1 U1109 ( .A1(n1662), .A2(n1567), .ZN(n1788) );
  OAI22_X1 U1106 ( .A1(B1[9]), .A2(n1432), .B1(B1[7]), .B2(n1661), .ZN(n1787)
         );
  AOI22_X1 U1104 ( .A1(n1783), .A2(n1784), .B1(n1785), .B2(n1786), .ZN(n1782)
         );
  XNOR2_X1 U1103 ( .A(n1752), .B(n1782), .ZN(n1754) );
  AOI221_X1 U1098 ( .B1(n1556), .B2(B1[3]), .C1(n1557), .C2(n1665), .A(n1780), 
        .ZN(n1749) );
  AOI22_X1 U1096 ( .A1(B1[0]), .A2(n1530), .B1(n1529), .B2(n1438), .ZN(n1778)
         );
  XNOR2_X1 U1100 ( .A(n1754), .B(n1753), .ZN(n1779) );
  XNOR2_X1 U1097 ( .A(n1779), .B(n1749), .ZN(n1751) );
  AOI22_X1 U1236 ( .A1(B1[0]), .A2(n1662), .B1(n1661), .B2(n1438), .ZN(n1866)
         );
  AOI221_X1 U1235 ( .B1(n1698), .B2(B1[1]), .C1(n1699), .C2(n1436), .A(n1866), 
        .ZN(n1525) );
  AOI22_X1 U1233 ( .A1(B1[3]), .A2(n1434), .B1(n1435), .B2(n1665), .ZN(n1865)
         );
  OAI21_X1 U1232 ( .B1(B1[2]), .B2(n1432), .A(n1865), .ZN(n1864) );
  AOI221_X1 U1248 ( .B1(n1698), .B2(B1[0]), .C1(n1699), .C2(n1438), .A(n1871), 
        .ZN(n1527) );
  OAI21_X1 U1240 ( .B1(B1[1]), .B2(n1432), .A(n1868), .ZN(n1867) );
  NOR2_X1 U1238 ( .A1(n1527), .A2(n1528), .ZN(p7_C[32]) );
  OAI221_X1 U863 ( .B1(B1[0]), .B2(n1437), .C1(n1438), .C2(n1439), .A(n1432), 
        .ZN(p7_final_product1[0]) );
  OAI221_X1 U1221 ( .B1(B1[1]), .B2(n1661), .C1(n1436), .C2(n1662), .A(n1861), 
        .ZN(n1520) );
  AOI22_X1 U1219 ( .A1(B1[4]), .A2(n1434), .B1(n1435), .B2(n1625), .ZN(n1860)
         );
  OAI21_X1 U1218 ( .B1(B1[3]), .B2(n1432), .A(n1860), .ZN(n1519) );
  XNOR2_X1 U1217 ( .A(n1520), .B(n1519), .ZN(n1522) );
  AOI22_X1 U1209 ( .A1(B1[1]), .A2(n1631), .B1(n1632), .B2(n1436), .ZN(n1857)
         );
  OAI221_X1 U1208 ( .B1(B1[0]), .B2(n1617), .C1(n1438), .C2(n1618), .A(n1857), 
        .ZN(n1515) );
  OAI21_X1 U1210 ( .B1(B1[4]), .B2(n1432), .A(n1858), .ZN(n1513) );
  NAND2_X1 U884 ( .A1(n1519), .A2(n1520), .ZN(n1518) );
  NAND2_X1 U1205 ( .A1(n1855), .A2(n1856), .ZN(p7_C[35]) );
  NAND2_X1 U882 ( .A1(n1513), .A2(n1514), .ZN(n1511) );
  AOI221_X1 U1198 ( .B1(n1438), .B2(n1598), .C1(B1[0]), .C2(n1597), .A(n1853), 
        .ZN(n1843) );
  OAI221_X1 U1196 ( .B1(B1[1]), .B2(n1617), .C1(n1436), .C2(n1618), .A(n1852), 
        .ZN(n1837) );
  OAI22_X1 U1180 ( .A1(B1[5]), .A2(n1432), .B1(B1[3]), .B2(n1661), .ZN(n1842)
         );
  AOI221_X1 U1179 ( .B1(n1434), .B2(B1[6]), .C1(n1435), .C2(n1591), .A(n1842), 
        .ZN(n1840) );
  AOI22_X1 U1178 ( .A1(B1[4]), .A2(n1698), .B1(n1699), .B2(n1625), .ZN(n1841)
         );
  OAI211_X1 U1177 ( .C1(n1662), .C2(n1665), .A(n1840), .B(n1841), .ZN(n1839)
         );
  OAI21_X1 U1176 ( .B1(n1837), .B2(n1838), .A(n1839), .ZN(n1505) );
  AOI22_X1 U1192 ( .A1(B1[0]), .A2(n1572), .B1(n1571), .B2(n1438), .ZN(n1848)
         );
  AOI221_X1 U1191 ( .B1(n1597), .B2(B1[1]), .C1(n1598), .C2(n1436), .A(n1848), 
        .ZN(n1507) );
  AOI22_X1 U1190 ( .A1(B1[4]), .A2(n1662), .B1(n1661), .B2(n1625), .ZN(n1847)
         );
  OAI22_X1 U1188 ( .A1(B1[6]), .A2(n1432), .B1(B1[7]), .B2(n1437), .ZN(n1846)
         );
  AOI21_X1 U1187 ( .B1(n1434), .B2(B1[7]), .A(n1846), .ZN(n1826) );
  XNOR2_X1 U1186 ( .A(n1825), .B(n1826), .ZN(n1844) );
  AOI221_X1 U1184 ( .B1(n1631), .B2(B1[3]), .C1(n1632), .C2(n1665), .A(n1845), 
        .ZN(n1827) );
  XNOR2_X1 U1183 ( .A(n1844), .B(n1827), .ZN(n1508) );
  OAI21_X1 U1195 ( .B1(reg2_reg[7]), .B2(n1512), .A(n1513), .ZN(n1850) );
  AOI222_X1 U1175 ( .A1(n1507), .A2(n1508), .B1(n1507), .B2(n1505), .C1(n1508), 
        .C2(n1505), .ZN(p7_C[37]) );
  AOI22_X1 U1174 ( .A1(B1[3]), .A2(n1618), .B1(n1617), .B2(n1665), .ZN(n1836)
         );
  AOI22_X1 U1172 ( .A1(B1[6]), .A2(n1698), .B1(n1699), .B2(n1591), .ZN(n1835)
         );
  OAI21_X1 U1168 ( .B1(B1[7]), .B2(n1432), .A(n1834), .ZN(n1820) );
  XNOR2_X1 U1167 ( .A(n1821), .B(n1820), .ZN(n1813) );
  XNOR2_X1 U1166 ( .A(n1833), .B(n1813), .ZN(n1814) );
  AOI22_X1 U1165 ( .A1(B1[1]), .A2(n1572), .B1(n1571), .B2(n1436), .ZN(n1832)
         );
  XNOR2_X1 U1156 ( .A(n1812), .B(n1809), .ZN(n1829) );
  AOI222_X1 U1153 ( .A1(n1825), .A2(n1826), .B1(n1825), .B2(n1827), .C1(n1826), 
        .C2(n1827), .ZN(n1824) );
  AOI22_X1 U1148 ( .A1(B1[4]), .A2(n1618), .B1(n1617), .B2(n1625), .ZN(n1822)
         );
  AOI22_X1 U1144 ( .A1(B1[7]), .A2(n1698), .B1(n1699), .B2(n1567), .ZN(n1819)
         );
  AOI22_X1 U1141 ( .A1(B1[9]), .A2(n1434), .B1(n1435), .B2(n1553), .ZN(n1818)
         );
  OAI21_X1 U1140 ( .B1(B1[8]), .B2(n1432), .A(n1818), .ZN(n1800) );
  AOI22_X1 U1138 ( .A1(B1[0]), .A2(n1547), .B1(n1546), .B2(n1438), .ZN(n1815)
         );
  AOI22_X1 U1135 ( .A1(B1[1]), .A2(n1547), .B1(n1546), .B2(n1436), .ZN(n1802)
         );
  AOI222_X1 U1118 ( .A1(n1497), .A2(n1498), .B1(n1497), .B2(n1495), .C1(n1498), 
        .C2(n1495), .ZN(p7_C[40]) );
  AOI222_X1 U1094 ( .A1(n1493), .A2(n1494), .B1(n1493), .B2(n1491), .C1(n1494), 
        .C2(n1491), .ZN(p7_C[41]) );
  AOI222_X1 U1045 ( .A1(n1485), .A2(n1486), .B1(n1485), .B2(n1483), .C1(n1486), 
        .C2(n1483), .ZN(p7_C[43]) );
  XNOR2_X1 U873 ( .A(n1471), .B(n1472), .ZN(p7_S[46]) );
  AOI222_X1 U1000 ( .A1(n1478), .A2(n1477), .B1(n1478), .B2(n1476), .C1(n1477), 
        .C2(n1476), .ZN(p7_C[45]) );
  XNOR2_X1 U871 ( .A(n1463), .B(n1464), .ZN(p7_S[48]) );
  AOI222_X1 U961 ( .A1(n1469), .A2(n1470), .B1(n1469), .B2(n1467), .C1(n1470), 
        .C2(n1467), .ZN(p7_C[47]) );
  XNOR2_X1 U869 ( .A(n1455), .B(n1456), .ZN(p7_S[50]) );
  AOI222_X1 U929 ( .A1(n1461), .A2(n1462), .B1(n1461), .B2(n1459), .C1(n1462), 
        .C2(n1459), .ZN(p7_C[49]) );
  XNOR2_X1 U867 ( .A(n1447), .B(n1448), .ZN(p7_S[52]) );
  AOI222_X1 U904 ( .A1(n1453), .A2(n1454), .B1(n1453), .B2(n1451), .C1(n1454), 
        .C2(n1451), .ZN(p7_C[51]) );
  XNOR2_X1 U864 ( .A(n1440), .B(n1441), .ZN(p7_S[54]) );
  AOI222_X1 U891 ( .A1(n1444), .A2(n1532), .B1(n1444), .B2(n1446), .C1(n1532), 
        .C2(n1446), .ZN(p7_C[53]) );
  NOR2_X1 U52 ( .A1(n1431), .A2(n1428), .ZN(n515) );
  NOR2_X1 U281 ( .A1(n3675), .A2(n3706), .ZN(n532) );
  OAI21_X1 U279 ( .B1(reg4_reg[11]), .B2(reg4_reg[12]), .A(n527), .ZN(n859) );
  AOI22_X1 U94 ( .A1(B3[11]), .A2(n527), .B1(n525), .B2(n635), .ZN(n634) );
  AOI221_X1 U93 ( .B1(n529), .B2(B3[12]), .C1(n530), .C2(n526), .A(n634), .ZN(
        n543) );
  OAI21_X1 U330 ( .B1(reg4_reg[9]), .B2(reg4_reg[10]), .A(n631), .ZN(n897) );
  AOI22_X1 U98 ( .A1(B3[13]), .A2(n639), .B1(n640), .B2(n531), .ZN(n632) );
  OAI221_X1 U97 ( .B1(B3[12]), .B2(n630), .C1(n526), .C2(n631), .A(n632), .ZN(
        n633) );
  OAI221_X1 U91 ( .B1(B3[13]), .B2(n630), .C1(n531), .C2(n631), .A(n632), .ZN(
        n542) );
  AOI22_X1 U64 ( .A1(B3[13]), .A2(n529), .B1(n530), .B2(n531), .ZN(n528) );
  OAI221_X1 U63 ( .B1(B3[12]), .B2(n525), .C1(n526), .C2(n527), .A(n528), .ZN(
        p9_final_product2_26_) );
  AOI221_X1 U115 ( .B1(n639), .B2(B3[11]), .C1(n640), .C2(n635), .A(n659), 
        .ZN(n653) );
  OAI21_X1 U366 ( .B1(reg4_reg[7]), .B2(reg4_reg[8]), .A(n648), .ZN(n932) );
  AOI22_X1 U114 ( .A1(B3[13]), .A2(n657), .B1(n658), .B2(n531), .ZN(n649) );
  OAI221_X1 U113 ( .B1(B3[12]), .B2(n647), .C1(n526), .C2(n648), .A(n649), 
        .ZN(n550) );
  XNOR2_X1 U109 ( .A(n651), .B(n652), .ZN(n552) );
  OAI21_X1 U407 ( .B1(reg4_reg[6]), .B2(reg4_reg[5]), .A(n673), .ZN(n955) );
  AOI22_X1 U144 ( .A1(B3[13]), .A2(n698), .B1(n699), .B2(n531), .ZN(n674) );
  OAI221_X1 U126 ( .B1(B3[13]), .B2(n672), .C1(n531), .C2(n673), .A(n674), 
        .ZN(n665) );
  AOI22_X1 U128 ( .A1(B3[11]), .A2(n648), .B1(n647), .B2(n635), .ZN(n675) );
  AOI221_X1 U127 ( .B1(n657), .B2(B3[12]), .C1(n658), .C2(n526), .A(n675), 
        .ZN(n671) );
  XNOR2_X1 U125 ( .A(n671), .B(n665), .ZN(n666) );
  XNOR2_X1 U122 ( .A(n666), .B(n664), .ZN(n667) );
  OAI221_X1 U143 ( .B1(B3[12]), .B2(n672), .C1(n526), .C2(n673), .A(n674), 
        .ZN(n662) );
  AOI22_X1 U117 ( .A1(n660), .A2(n661), .B1(n662), .B2(n663), .ZN(n555) );
  XNOR2_X1 U72 ( .A(n552), .B(n553), .ZN(p9_S[51]) );
  AOI22_X1 U163 ( .A1(B3[11]), .A2(n673), .B1(n672), .B2(n635), .ZN(n721) );
  AOI221_X1 U162 ( .B1(n698), .B2(B3[12]), .C1(n699), .C2(n526), .A(n721), 
        .ZN(n700) );
  OAI21_X1 U432 ( .B1(reg4_reg[3]), .B2(reg4_reg[4]), .A(n719), .ZN(n964) );
  AOI22_X1 U177 ( .A1(B3[13]), .A2(n732), .B1(n733), .B2(n531), .ZN(n720) );
  OAI221_X1 U161 ( .B1(B3[13]), .B2(n718), .C1(n531), .C2(n719), .A(n720), 
        .ZN(n701) );
  XNOR2_X1 U160 ( .A(n700), .B(n701), .ZN(n702) );
  OAI22_X1 U145 ( .A1(n700), .A2(n701), .B1(n702), .B2(n703), .ZN(n682) );
  AOI221_X1 U141 ( .B1(n657), .B2(B3[11]), .C1(n658), .C2(n635), .A(n697), 
        .ZN(n684) );
  AOI22_X1 U130 ( .A1(n680), .A2(n681), .B1(n682), .B2(n683), .ZN(n558) );
  OAI221_X1 U135 ( .B1(B3[6]), .B2(n525), .C1(n692), .C2(n527), .A(n693), .ZN(
        n677) );
  AOI22_X1 U129 ( .A1(n676), .A2(n677), .B1(n678), .B2(n679), .ZN(n559) );
  AOI222_X1 U119 ( .A1(n558), .A2(n559), .B1(n558), .B2(n556), .C1(n559), .C2(
        n556), .ZN(p9_C[50]) );
  OAI21_X1 U458 ( .B1(reg4_reg[1]), .B2(reg4_reg[2]), .A(n763), .ZN(n973) );
  NAND2_X1 U454 ( .A1(reg4_reg[3]), .A2(n973), .ZN(n762) );
  AOI22_X1 U227 ( .A1(B3[13]), .A2(n799), .B1(n800), .B2(n531), .ZN(n764) );
  OAI221_X1 U197 ( .B1(B3[13]), .B2(n762), .C1(n531), .C2(n763), .A(n764), 
        .ZN(n738) );
  AOI22_X1 U196 ( .A1(B3[12]), .A2(n732), .B1(n733), .B2(n526), .ZN(n761) );
  OAI221_X1 U195 ( .B1(B3[11]), .B2(n718), .C1(n635), .C2(n719), .A(n761), 
        .ZN(n760) );
  AOI22_X1 U192 ( .A1(B3[6]), .A2(n639), .B1(n640), .B2(n692), .ZN(n757) );
  AOI22_X1 U182 ( .A1(n739), .A2(n740), .B1(n741), .B2(n742), .ZN(n708) );
  NAND2_X1 U181 ( .A1(n735), .A2(n738), .ZN(n737) );
  OAI21_X1 U180 ( .B1(n735), .B2(n736), .A(n737), .ZN(n729) );
  AOI221_X1 U178 ( .B1(n698), .B2(B3[11]), .C1(n699), .C2(n635), .A(n734), 
        .ZN(n722) );
  OAI221_X1 U176 ( .B1(B3[12]), .B2(n718), .C1(n526), .C2(n719), .A(n720), 
        .ZN(n686) );
  XNOR2_X1 U175 ( .A(n722), .B(n686), .ZN(n723) );
  AOI22_X1 U171 ( .A1(B3[6]), .A2(n631), .B1(n630), .B2(n692), .ZN(n728) );
  XNOR2_X1 U169 ( .A(n727), .B(n705), .ZN(n706) );
  AOI22_X1 U168 ( .A1(B3[4]), .A2(n527), .B1(n525), .B2(n726), .ZN(n725) );
  XNOR2_X1 U166 ( .A(n706), .B(n704), .ZN(n568) );
  OAI221_X1 U226 ( .B1(B3[12]), .B2(n762), .C1(n526), .C2(n763), .A(n764), 
        .ZN(n746) );
  AOI221_X1 U228 ( .B1(n732), .B2(B3[11]), .C1(n733), .C2(n635), .A(n801), 
        .ZN(n798) );
  XNOR2_X1 U225 ( .A(n798), .B(n746), .ZN(n756) );
  AOI22_X1 U218 ( .A1(B3[4]), .A2(n631), .B1(n630), .B2(n726), .ZN(n794) );
  AOI22_X1 U224 ( .A1(B3[6]), .A2(n648), .B1(n647), .B2(n692), .ZN(n797) );
  XNOR2_X1 U222 ( .A(n756), .B(n769), .ZN(n795) );
  XNOR2_X1 U219 ( .A(n795), .B(n755), .ZN(n770) );
  AOI22_X1 U186 ( .A1(n748), .A2(n749), .B1(n750), .B2(n751), .ZN(n570) );
  AOI22_X1 U201 ( .A1(B3[4]), .A2(n529), .B1(n530), .B2(n726), .ZN(n767) );
  OAI221_X1 U200 ( .B1(B3[3]), .B2(n525), .C1(n766), .C2(n527), .A(n767), .ZN(
        n745) );
  AOI22_X1 U185 ( .A1(n744), .A2(n745), .B1(n746), .B2(n747), .ZN(n571) );
  XNOR2_X1 U76 ( .A(n568), .B(n569), .ZN(p9_S[47]) );
  XNOR2_X1 U216 ( .A(n770), .B(n768), .ZN(n776) );
  NAND2_X1 U450 ( .A1(n3701), .A2(reg4_reg[0]), .ZN(n540) );
  AOI22_X1 U241 ( .A1(B3[13]), .A2(n535), .B1(reg4_reg[1]), .B2(n531), .ZN(
        n802) );
  AOI22_X1 U239 ( .A1(B3[11]), .A2(n763), .B1(n762), .B2(n635), .ZN(n821) );
  AOI221_X1 U238 ( .B1(n799), .B2(B3[12]), .C1(n800), .C2(n526), .A(n821), 
        .ZN(n820) );
  AOI22_X1 U235 ( .A1(B3[6]), .A2(n657), .B1(n658), .B2(n692), .ZN(n817) );
  OAI22_X1 U230 ( .A1(n802), .A2(n803), .B1(n804), .B2(n805), .ZN(n793) );
  AOI22_X1 U248 ( .A1(B3[3]), .A2(n631), .B1(n630), .B2(n766), .ZN(n824) );
  AOI22_X1 U246 ( .A1(B3[1]), .A2(n527), .B1(n525), .B2(n537), .ZN(n823) );
  NOR2_X1 U215 ( .A1(n774), .A2(n775), .ZN(n792) );
  XNOR2_X1 U214 ( .A(n778), .B(n792), .ZN(n786) );
  XNOR2_X1 U210 ( .A(n786), .B(n777), .ZN(n771) );
  AOI22_X1 U209 ( .A1(B3[3]), .A2(n529), .B1(n530), .B2(n766), .ZN(n785) );
  OAI21_X1 U203 ( .B1(n774), .B2(n775), .A(n771), .ZN(n773) );
  OAI21_X1 U202 ( .B1(n771), .B2(n772), .A(n773), .ZN(n575) );
  AOI222_X1 U189 ( .A1(n574), .A2(n575), .B1(n574), .B2(n572), .C1(n575), .C2(
        n572), .ZN(p9_C[46]) );
  AOI22_X1 U440 ( .A1(B3[0]), .A2(n763), .B1(n762), .B2(n539), .ZN(n967) );
  AOI221_X1 U439 ( .B1(n799), .B2(B3[1]), .C1(n800), .C2(n537), .A(n967), .ZN(
        n626) );
  NAND2_X1 U451 ( .A1(reg4_reg[1]), .A2(n3705), .ZN(n533) );
  NAND2_X1 U448 ( .A1(reg4_reg[0]), .A2(reg4_reg[1]), .ZN(n538) );
  AOI22_X1 U437 ( .A1(B3[3]), .A2(n535), .B1(n536), .B2(n766), .ZN(n966) );
  OAI21_X1 U436 ( .B1(B3[2]), .B2(n533), .A(n966), .ZN(n965) );
  AOI221_X1 U452 ( .B1(n799), .B2(B3[0]), .C1(n800), .C2(n539), .A(n972), .ZN(
        n628) );
  OAI21_X1 U444 ( .B1(B3[1]), .B2(n533), .A(n969), .ZN(n968) );
  NOR2_X1 U442 ( .A1(n628), .A2(n629), .ZN(p9_C[32]) );
  OAI221_X1 U425 ( .B1(B3[1]), .B2(n762), .C1(n537), .C2(n763), .A(n962), .ZN(
        n621) );
  AOI22_X1 U423 ( .A1(B3[4]), .A2(n535), .B1(n536), .B2(n726), .ZN(n961) );
  OAI21_X1 U422 ( .B1(B3[3]), .B2(n533), .A(n961), .ZN(n620) );
  XNOR2_X1 U421 ( .A(n621), .B(n620), .ZN(n623) );
  XNOR2_X1 U89 ( .A(n622), .B(n623), .ZN(p9_S[34]) );
  NOR2_X1 U434 ( .A1(n626), .A2(n627), .ZN(p9_C[33]) );
  AOI22_X1 U413 ( .A1(B3[1]), .A2(n732), .B1(n733), .B2(n537), .ZN(n958) );
  OAI221_X1 U412 ( .B1(B3[0]), .B2(n718), .C1(n539), .C2(n719), .A(n958), .ZN(
        n616) );
  AOI221_X1 U418 ( .B1(n799), .B2(B3[3]), .C1(n800), .C2(n766), .A(n960), .ZN(
        n950) );
  OAI21_X1 U414 ( .B1(B3[4]), .B2(n533), .A(n959), .ZN(n614) );
  NAND2_X1 U88 ( .A1(n620), .A2(n621), .ZN(n619) );
  NAND2_X1 U409 ( .A1(n956), .A2(n957), .ZN(p9_C[35]) );
  NAND2_X1 U86 ( .A1(n614), .A2(n615), .ZN(n612) );
  AOI221_X1 U402 ( .B1(n539), .B2(n699), .C1(B3[0]), .C2(n698), .A(n954), .ZN(
        n944) );
  OAI221_X1 U400 ( .B1(B3[1]), .B2(n718), .C1(n537), .C2(n719), .A(n953), .ZN(
        n938) );
  OAI22_X1 U384 ( .A1(B3[5]), .A2(n533), .B1(B3[3]), .B2(n762), .ZN(n943) );
  AOI221_X1 U383 ( .B1(n535), .B2(B3[6]), .C1(n536), .C2(n692), .A(n943), .ZN(
        n941) );
  AOI22_X1 U382 ( .A1(B3[4]), .A2(n799), .B1(n800), .B2(n726), .ZN(n942) );
  OAI211_X1 U381 ( .C1(n763), .C2(n766), .A(n941), .B(n942), .ZN(n940) );
  OAI21_X1 U380 ( .B1(n938), .B2(n939), .A(n940), .ZN(n606) );
  AOI22_X1 U396 ( .A1(B3[0]), .A2(n673), .B1(n672), .B2(n539), .ZN(n949) );
  AOI221_X1 U395 ( .B1(n698), .B2(B3[1]), .C1(n699), .C2(n537), .A(n949), .ZN(
        n608) );
  AOI22_X1 U394 ( .A1(B3[4]), .A2(n763), .B1(n762), .B2(n726), .ZN(n948) );
  OAI22_X1 U392 ( .A1(B3[6]), .A2(n533), .B1(B3[7]), .B2(n538), .ZN(n947) );
  AOI21_X1 U391 ( .B1(n535), .B2(B3[7]), .A(n947), .ZN(n927) );
  XNOR2_X1 U390 ( .A(n926), .B(n927), .ZN(n945) );
  AOI221_X1 U388 ( .B1(n732), .B2(B3[3]), .C1(n733), .C2(n766), .A(n946), .ZN(
        n928) );
  XNOR2_X1 U387 ( .A(n945), .B(n928), .ZN(n609) );
  OAI21_X1 U399 ( .B1(reg4_reg[7]), .B2(n613), .A(n614), .ZN(n951) );
  OAI22_X1 U397 ( .A1(n950), .A2(n951), .B1(n952), .B2(n3697), .ZN(p9_C[36])
         );
  AOI222_X1 U379 ( .A1(n608), .A2(n609), .B1(n608), .B2(n606), .C1(n609), .C2(
        n606), .ZN(p9_C[37]) );
  AOI22_X1 U378 ( .A1(B3[3]), .A2(n719), .B1(n718), .B2(n766), .ZN(n937) );
  OAI21_X1 U372 ( .B1(B3[7]), .B2(n533), .A(n935), .ZN(n921) );
  XNOR2_X1 U370 ( .A(n934), .B(n914), .ZN(n915) );
  AOI22_X1 U369 ( .A1(B3[1]), .A2(n673), .B1(n672), .B2(n537), .ZN(n933) );
  XNOR2_X1 U360 ( .A(n913), .B(n910), .ZN(n930) );
  AOI222_X1 U357 ( .A1(n926), .A2(n927), .B1(n926), .B2(n928), .C1(n927), .C2(
        n928), .ZN(n925) );
  AOI22_X1 U352 ( .A1(B3[4]), .A2(n719), .B1(n718), .B2(n726), .ZN(n923) );
  OAI21_X1 U344 ( .B1(B3[8]), .B2(n533), .A(n919), .ZN(n901) );
  AOI22_X1 U342 ( .A1(B3[0]), .A2(n648), .B1(n647), .B2(n539), .ZN(n916) );
  NOR2_X1 U355 ( .A1(n605), .A2(n604), .ZN(p9_C[38]) );
  AOI22_X1 U339 ( .A1(B3[1]), .A2(n648), .B1(n647), .B2(n537), .ZN(n903) );
  AOI22_X1 U336 ( .A1(B3[3]), .A2(n673), .B1(n672), .B2(n766), .ZN(n900) );
  AOI221_X1 U320 ( .B1(n799), .B2(B3[9]), .C1(n800), .C2(n654), .A(n893), .ZN(
        n870) );
  OAI22_X1 U319 ( .A1(B3[11]), .A2(n538), .B1(B3[10]), .B2(n533), .ZN(n892) );
  AOI21_X1 U318 ( .B1(B3[11]), .B2(n535), .A(n892), .ZN(n871) );
  XNOR2_X1 U314 ( .A(n890), .B(n872), .ZN(n853) );
  OAI22_X1 U310 ( .A1(B3[9]), .A2(n533), .B1(B3[7]), .B2(n762), .ZN(n888) );
  XNOR2_X1 U307 ( .A(n853), .B(n883), .ZN(n855) );
  AOI22_X1 U306 ( .A1(B3[4]), .A2(n673), .B1(n672), .B2(n726), .ZN(n882) );
  XNOR2_X1 U304 ( .A(n855), .B(n854), .ZN(n880) );
  AOI221_X1 U302 ( .B1(n657), .B2(B3[3]), .C1(n658), .C2(n766), .A(n881), .ZN(
        n850) );
  XNOR2_X1 U301 ( .A(n880), .B(n850), .ZN(n852) );
  AOI22_X1 U300 ( .A1(B3[0]), .A2(n631), .B1(n630), .B2(n539), .ZN(n879) );
  AOI22_X1 U297 ( .A1(B3[1]), .A2(n631), .B1(n630), .B2(n537), .ZN(n873) );
  OAI22_X1 U294 ( .A1(B3[11]), .A2(n533), .B1(B3[12]), .B2(n538), .ZN(n869) );
  AOI21_X1 U293 ( .B1(B3[12]), .B2(n535), .A(n869), .ZN(n831) );
  AOI22_X1 U283 ( .A1(B3[3]), .A2(n648), .B1(n647), .B2(n766), .ZN(n863) );
  XNOR2_X1 U267 ( .A(n810), .B(n807), .ZN(n829) );
  OAI221_X1 U265 ( .B1(B3[6]), .B2(n672), .C1(n692), .C2(n673), .A(n840), .ZN(
        n813) );
  AOI221_X1 U262 ( .B1(n799), .B2(B3[11]), .C1(n800), .C2(n635), .A(n839), 
        .ZN(n837) );
  AOI22_X1 U260 ( .A1(B3[13]), .A2(n535), .B1(n536), .B2(n531), .ZN(n838) );
  OAI21_X1 U259 ( .B1(B3[12]), .B2(n533), .A(n838), .ZN(n825) );
  XNOR2_X1 U258 ( .A(n837), .B(n825), .ZN(n827) );
  OAI221_X1 U254 ( .B1(B3[4]), .B2(n647), .C1(n726), .C2(n648), .A(n834), .ZN(
        n814) );
  XNOR2_X1 U253 ( .A(n815), .B(n814), .ZN(n809) );
  AOI22_X1 U252 ( .A1(B3[0]), .A2(n527), .B1(n525), .B2(n539), .ZN(n828) );
  XNOR2_X1 U250 ( .A(n808), .B(n806), .ZN(n584) );
  XNOR2_X1 U80 ( .A(n584), .B(n585), .ZN(p9_S[43]) );
  XNOR2_X1 U244 ( .A(n774), .B(n775), .ZN(n816) );
  AOI222_X1 U249 ( .A1(n586), .A2(n587), .B1(n586), .B2(n584), .C1(n587), .C2(
        n584), .ZN(p9_C[43]) );
  XNOR2_X1 U78 ( .A(n578), .B(n579), .ZN(n576) );
  XNOR2_X1 U77 ( .A(n572), .B(n573), .ZN(p9_S[46]) );
  AOI222_X1 U204 ( .A1(n579), .A2(n578), .B1(n579), .B2(n577), .C1(n578), .C2(
        n577), .ZN(p9_C[45]) );
  OAI22_X1 U164 ( .A1(n722), .A2(n686), .B1(n723), .B2(n724), .ZN(n716) );
  XNOR2_X1 U157 ( .A(n702), .B(n703), .ZN(n689) );
  XNOR2_X1 U156 ( .A(n716), .B(n689), .ZN(n691) );
  XNOR2_X1 U153 ( .A(n691), .B(n690), .ZN(n711) );
  AOI22_X1 U147 ( .A1(n707), .A2(n708), .B1(n709), .B2(n710), .ZN(n567) );
  XNOR2_X1 U75 ( .A(n564), .B(n565), .ZN(p9_S[48]) );
  AOI222_X1 U165 ( .A1(n570), .A2(n571), .B1(n570), .B2(n568), .C1(n571), .C2(
        n568), .ZN(p9_C[47]) );
  AOI22_X1 U134 ( .A1(n685), .A2(n686), .B1(n687), .B2(n688), .ZN(n560) );
  XNOR2_X1 U74 ( .A(n560), .B(n561), .ZN(p9_S[49]) );
  AOI222_X1 U146 ( .A1(n566), .A2(n567), .B1(n566), .B2(n564), .C1(n567), .C2(
        n564), .ZN(p9_C[48]) );
  XNOR2_X1 U73 ( .A(n556), .B(n557), .ZN(p9_S[50]) );
  AOI222_X1 U133 ( .A1(n562), .A2(n563), .B1(n562), .B2(n560), .C1(n563), .C2(
        n560), .ZN(p9_C[49]) );
  OAI22_X1 U107 ( .A1(n651), .A2(n652), .B1(n653), .B2(n550), .ZN(n551) );
  AOI22_X1 U105 ( .A1(B3[12]), .A2(n639), .B1(n640), .B2(n526), .ZN(n650) );
  OAI221_X1 U104 ( .B1(B3[11]), .B2(n630), .C1(n635), .C2(n631), .A(n650), 
        .ZN(n637) );
  OAI221_X1 U103 ( .B1(B3[13]), .B2(n647), .C1(n531), .C2(n648), .A(n649), 
        .ZN(n646) );
  XNOR2_X1 U71 ( .A(n548), .B(n549), .ZN(p9_S[52]) );
  AOI222_X1 U108 ( .A1(n554), .A2(n555), .B1(n554), .B2(n552), .C1(n555), .C2(
        n552), .ZN(p9_C[51]) );
  AOI221_X1 U99 ( .B1(n529), .B2(B3[11]), .C1(n530), .C2(n635), .A(n641), .ZN(
        n545) );
  AOI22_X1 U96 ( .A1(n636), .A2(n637), .B1(reg4_reg[13]), .B2(n638), .ZN(n547)
         );
  XNOR2_X1 U70 ( .A(n544), .B(n547), .ZN(n546) );
  XNOR2_X1 U69 ( .A(n545), .B(n546), .ZN(p9_S[53]) );
  AOI222_X1 U101 ( .A1(n643), .A2(n644), .B1(n643), .B2(n549), .C1(n644), .C2(
        n549), .ZN(p9_C[52]) );
  XNOR2_X1 U68 ( .A(n541), .B(n542), .ZN(p9_S[54]) );
  AOI222_X1 U95 ( .A1(n545), .A2(n633), .B1(n545), .B2(n547), .C1(n633), .C2(
        n547), .ZN(p9_C[53]) );
  NOR2_X1 U56 ( .A1(n532), .A2(n529), .ZN(n519) );
  OAI21_X1 U678 ( .B1(reg3_reg[11]), .B2(reg3_reg[12]), .A(n977), .ZN(n1309)
         );
  AOI22_X1 U493 ( .A1(B2[11]), .A2(n977), .B1(n975), .B2(n1085), .ZN(n1084) );
  AOI221_X1 U492 ( .B1(n979), .B2(B2[12]), .C1(n980), .C2(n976), .A(n1084), 
        .ZN(n993) );
  OAI21_X1 U728 ( .B1(reg3_reg[9]), .B2(reg3_reg[10]), .A(n1081), .ZN(n1346)
         );
  AOI22_X1 U497 ( .A1(B2[13]), .A2(n1089), .B1(n1090), .B2(n981), .ZN(n1082)
         );
  OAI221_X1 U496 ( .B1(B2[12]), .B2(n1080), .C1(n976), .C2(n1081), .A(n1082), 
        .ZN(n1083) );
  OAI221_X1 U490 ( .B1(B2[13]), .B2(n1080), .C1(n981), .C2(n1081), .A(n1082), 
        .ZN(n992) );
  AOI222_X1 U489 ( .A1(n993), .A2(n994), .B1(n993), .B2(n992), .C1(n994), .C2(
        n992), .ZN(p8_C[54]) );
  AOI22_X1 U523 ( .A1(B2[9]), .A2(n1081), .B1(n1080), .B2(n1104), .ZN(n1120)
         );
  OAI21_X1 U805 ( .B1(reg3_reg[6]), .B2(reg3_reg[5]), .A(n1123), .ZN(n1404) );
  AOI22_X1 U543 ( .A1(B2[13]), .A2(n1148), .B1(n1149), .B2(n981), .ZN(n1124)
         );
  OAI221_X1 U525 ( .B1(B2[13]), .B2(n1122), .C1(n981), .C2(n1123), .A(n1124), 
        .ZN(n1115) );
  OAI21_X1 U764 ( .B1(reg3_reg[7]), .B2(reg3_reg[8]), .A(n1098), .ZN(n1381) );
  AOI22_X1 U527 ( .A1(B2[11]), .A2(n1098), .B1(n1097), .B2(n1085), .ZN(n1125)
         );
  AOI221_X1 U526 ( .B1(n1107), .B2(B2[12]), .C1(n1108), .C2(n976), .A(n1125), 
        .ZN(n1121) );
  XNOR2_X1 U524 ( .A(n1121), .B(n1115), .ZN(n1116) );
  XNOR2_X1 U521 ( .A(n1116), .B(n1114), .ZN(n1117) );
  OAI221_X1 U519 ( .B1(B2[7]), .B2(n975), .C1(n1118), .C2(n977), .A(n1119), 
        .ZN(n1111) );
  OAI221_X1 U542 ( .B1(B2[12]), .B2(n1122), .C1(n976), .C2(n1123), .A(n1124), 
        .ZN(n1112) );
  AOI22_X1 U516 ( .A1(n1110), .A2(n1111), .B1(n1112), .B2(n1113), .ZN(n1005)
         );
  AOI221_X1 U514 ( .B1(n1089), .B2(B2[11]), .C1(n1090), .C2(n1085), .A(n1109), 
        .ZN(n1103) );
  AOI22_X1 U513 ( .A1(B2[13]), .A2(n1107), .B1(n1108), .B2(n981), .ZN(n1099)
         );
  OAI221_X1 U512 ( .B1(B2[12]), .B2(n1097), .C1(n976), .C2(n1098), .A(n1099), 
        .ZN(n1000) );
  AOI221_X1 U509 ( .B1(n979), .B2(B2[9]), .C1(n980), .C2(n1104), .A(n1105), 
        .ZN(n1102) );
  XNOR2_X1 U508 ( .A(n1101), .B(n1102), .ZN(n1002) );
  AOI222_X1 U507 ( .A1(n1004), .A2(n1005), .B1(n1004), .B2(n1002), .C1(n1005), 
        .C2(n1002), .ZN(p8_C[51]) );
  OAI22_X1 U506 ( .A1(n1101), .A2(n1102), .B1(n1103), .B2(n1000), .ZN(n1001)
         );
  AOI22_X1 U504 ( .A1(B2[12]), .A2(n1089), .B1(n1090), .B2(n976), .ZN(n1100)
         );
  OAI221_X1 U503 ( .B1(B2[11]), .B2(n1080), .C1(n1085), .C2(n1081), .A(n1100), 
        .ZN(n1087) );
  OAI221_X1 U502 ( .B1(B2[13]), .B2(n1097), .C1(n981), .C2(n1098), .A(n1099), 
        .ZN(n1096) );
  XNOR2_X1 U470 ( .A(n998), .B(n999), .ZN(p8_S[52]) );
  XNOR2_X1 U471 ( .A(n1002), .B(n1003), .ZN(p8_S[51]) );
  AOI22_X1 U562 ( .A1(B2[11]), .A2(n1123), .B1(n1122), .B2(n1085), .ZN(n1171)
         );
  AOI221_X1 U561 ( .B1(n1148), .B2(B2[12]), .C1(n1149), .C2(n976), .A(n1171), 
        .ZN(n1150) );
  OAI21_X1 U830 ( .B1(reg3_reg[3]), .B2(reg3_reg[4]), .A(n1169), .ZN(n1413) );
  AOI22_X1 U576 ( .A1(B2[13]), .A2(n1182), .B1(n1183), .B2(n981), .ZN(n1170)
         );
  OAI221_X1 U560 ( .B1(B2[13]), .B2(n1168), .C1(n981), .C2(n1169), .A(n1170), 
        .ZN(n1151) );
  XNOR2_X1 U559 ( .A(n1150), .B(n1151), .ZN(n1152) );
  AOI22_X1 U558 ( .A1(B2[9]), .A2(n1098), .B1(n1097), .B2(n1104), .ZN(n1167)
         );
  OAI22_X1 U544 ( .A1(n1150), .A2(n1151), .B1(n1152), .B2(n1153), .ZN(n1132)
         );
  AOI221_X1 U540 ( .B1(n1107), .B2(B2[11]), .C1(n1108), .C2(n1085), .A(n1147), 
        .ZN(n1134) );
  AOI22_X1 U529 ( .A1(n1130), .A2(n1131), .B1(n1132), .B2(n1133), .ZN(n1008)
         );
  AOI221_X1 U538 ( .B1(n1089), .B2(B2[9]), .C1(n1090), .C2(n1104), .A(n1146), 
        .ZN(n1145) );
  AOI22_X1 U535 ( .A1(B2[7]), .A2(n979), .B1(n980), .B2(n1118), .ZN(n1143) );
  OAI221_X1 U534 ( .B1(B2[6]), .B2(n975), .C1(n1142), .C2(n977), .A(n1143), 
        .ZN(n1127) );
  AOI22_X1 U528 ( .A1(n1126), .A2(n1127), .B1(n1128), .B2(n1129), .ZN(n1009)
         );
  AOI221_X1 U577 ( .B1(n1148), .B2(B2[11]), .C1(n1149), .C2(n1085), .A(n1184), 
        .ZN(n1172) );
  OAI221_X1 U575 ( .B1(B2[12]), .B2(n1168), .C1(n976), .C2(n1169), .A(n1170), 
        .ZN(n1136) );
  XNOR2_X1 U574 ( .A(n1172), .B(n1136), .ZN(n1173) );
  AOI22_X1 U573 ( .A1(B2[9]), .A2(n1107), .B1(n1108), .B2(n1104), .ZN(n1181)
         );
  OAI22_X1 U563 ( .A1(n1172), .A2(n1136), .B1(n1173), .B2(n1174), .ZN(n1166)
         );
  XNOR2_X1 U556 ( .A(n1152), .B(n1153), .ZN(n1139) );
  XNOR2_X1 U555 ( .A(n1166), .B(n1139), .ZN(n1141) );
  AOI22_X1 U554 ( .A1(B2[7]), .A2(n1081), .B1(n1080), .B2(n1118), .ZN(n1165)
         );
  XNOR2_X1 U552 ( .A(n1141), .B(n1140), .ZN(n1161) );
  AOI22_X1 U533 ( .A1(n1135), .A2(n1136), .B1(n1137), .B2(n1138), .ZN(n1010)
         );
  XNOR2_X1 U473 ( .A(n1010), .B(n1011), .ZN(p8_S[49]) );
  OAI21_X1 U856 ( .B1(reg3_reg[1]), .B2(reg3_reg[2]), .A(n1213), .ZN(n1422) );
  NAND2_X1 U852 ( .A1(reg3_reg[3]), .A2(n1422), .ZN(n1212) );
  AOI22_X1 U626 ( .A1(B2[13]), .A2(n1249), .B1(n1250), .B2(n981), .ZN(n1214)
         );
  OAI221_X1 U596 ( .B1(B2[13]), .B2(n1212), .C1(n981), .C2(n1213), .A(n1214), 
        .ZN(n1188) );
  AOI22_X1 U595 ( .A1(B2[12]), .A2(n1182), .B1(n1183), .B2(n976), .ZN(n1211)
         );
  OAI221_X1 U594 ( .B1(B2[11]), .B2(n1168), .C1(n1085), .C2(n1169), .A(n1211), 
        .ZN(n1210) );
  OAI221_X1 U592 ( .B1(B2[9]), .B2(n1122), .C1(n1104), .C2(n1123), .A(n1209), 
        .ZN(n1186) );
  NAND2_X1 U580 ( .A1(n1185), .A2(n1188), .ZN(n1187) );
  OAI21_X1 U579 ( .B1(n1185), .B2(n1186), .A(n1187), .ZN(n1179) );
  AOI22_X1 U598 ( .A1(B2[7]), .A2(n1098), .B1(n1097), .B2(n1118), .ZN(n1215)
         );
  AOI22_X1 U591 ( .A1(B2[6]), .A2(n1089), .B1(n1090), .B2(n1142), .ZN(n1207)
         );
  AOI22_X1 U581 ( .A1(n1189), .A2(n1190), .B1(n1191), .B2(n1192), .ZN(n1158)
         );
  AOI22_X1 U546 ( .A1(n1157), .A2(n1158), .B1(n1159), .B2(n1160), .ZN(n1017)
         );
  AOI22_X1 U567 ( .A1(B2[4]), .A2(n977), .B1(n975), .B2(n1176), .ZN(n1175) );
  AOI22_X1 U570 ( .A1(B2[6]), .A2(n1081), .B1(n1080), .B2(n1142), .ZN(n1178)
         );
  AOI221_X1 U569 ( .B1(n1089), .B2(B2[7]), .C1(n1090), .C2(n1118), .A(n1178), 
        .ZN(n1155) );
  XNOR2_X1 U568 ( .A(n1177), .B(n1155), .ZN(n1156) );
  AOI222_X1 U545 ( .A1(n1016), .A2(n1017), .B1(n1016), .B2(n1014), .C1(n1017), 
        .C2(n1014), .ZN(p8_C[48]) );
  XNOR2_X1 U565 ( .A(n1156), .B(n1154), .ZN(n1018) );
  AOI221_X1 U619 ( .B1(n1148), .B2(B2[9]), .C1(n1149), .C2(n1104), .A(n1246), 
        .ZN(n1205) );
  OAI221_X1 U625 ( .B1(B2[12]), .B2(n1212), .C1(n976), .C2(n1213), .A(n1214), 
        .ZN(n1196) );
  AOI221_X1 U627 ( .B1(n1182), .B2(B2[11]), .C1(n1183), .C2(n1085), .A(n1251), 
        .ZN(n1248) );
  XNOR2_X1 U624 ( .A(n1248), .B(n1196), .ZN(n1206) );
  AOI22_X1 U617 ( .A1(B2[4]), .A2(n1081), .B1(n1080), .B2(n1176), .ZN(n1244)
         );
  AOI22_X1 U623 ( .A1(B2[6]), .A2(n1098), .B1(n1097), .B2(n1142), .ZN(n1247)
         );
  XNOR2_X1 U621 ( .A(n1206), .B(n1219), .ZN(n1245) );
  XNOR2_X1 U618 ( .A(n1245), .B(n1205), .ZN(n1220) );
  AOI22_X1 U585 ( .A1(n1198), .A2(n1199), .B1(n1200), .B2(n1201), .ZN(n1020)
         );
  AOI22_X1 U600 ( .A1(B2[4]), .A2(n979), .B1(n980), .B2(n1176), .ZN(n1217) );
  OAI221_X1 U599 ( .B1(B2[3]), .B2(n975), .C1(n3827), .C2(n977), .A(n1217), 
        .ZN(n1195) );
  AOI22_X1 U584 ( .A1(n1194), .A2(n1195), .B1(n1196), .B2(n1197), .ZN(n1021)
         );
  XNOR2_X1 U475 ( .A(n1018), .B(n1019), .ZN(p8_S[47]) );
  XNOR2_X1 U615 ( .A(n1220), .B(n1218), .ZN(n1226) );
  AOI221_X1 U641 ( .B1(n1148), .B2(B2[8]), .C1(n1149), .C2(n1106), .A(n1272), 
        .ZN(n1241) );
  NAND2_X1 U848 ( .A1(n3700), .A2(reg3_reg[0]), .ZN(n990) );
  AOI22_X1 U640 ( .A1(B2[13]), .A2(n985), .B1(reg3_reg[1]), .B2(n981), .ZN(
        n1252) );
  AOI22_X1 U638 ( .A1(B2[11]), .A2(n1213), .B1(n1212), .B2(n1085), .ZN(n1271)
         );
  AOI221_X1 U637 ( .B1(n1249), .B2(B2[12]), .C1(n1250), .C2(n976), .A(n1271), 
        .ZN(n1270) );
  AOI22_X1 U634 ( .A1(B2[6]), .A2(n1107), .B1(n1108), .B2(n1142), .ZN(n1267)
         );
  AOI22_X1 U647 ( .A1(B2[3]), .A2(n1081), .B1(n1080), .B2(n3827), .ZN(n1274)
         );
  AOI22_X1 U645 ( .A1(B2[1]), .A2(n977), .B1(n975), .B2(n987), .ZN(n1273) );
  NOR2_X1 U614 ( .A1(n1224), .A2(n1225), .ZN(n1242) );
  XNOR2_X1 U613 ( .A(n1228), .B(n1242), .ZN(n1236) );
  XNOR2_X1 U609 ( .A(n1236), .B(n1227), .ZN(n1221) );
  AOI22_X1 U608 ( .A1(B2[3]), .A2(n979), .B1(n980), .B2(n3827), .ZN(n1235) );
  OAI21_X1 U602 ( .B1(n1224), .B2(n1225), .A(n1221), .ZN(n1223) );
  OAI21_X1 U601 ( .B1(n1221), .B2(n1222), .A(n1223), .ZN(n1025) );
  AOI222_X1 U588 ( .A1(n1024), .A2(n1025), .B1(n1024), .B2(n1022), .C1(n1025), 
        .C2(n1022), .ZN(p8_C[46]) );
  AOI22_X1 U665 ( .A1(B2[7]), .A2(n1148), .B1(n1149), .B2(n1118), .ZN(n1290)
         );
  OAI221_X1 U664 ( .B1(B2[6]), .B2(n1122), .C1(n1142), .C2(n1123), .A(n1290), 
        .ZN(n1263) );
  OAI221_X1 U653 ( .B1(B2[4]), .B2(n1097), .C1(n1176), .C2(n1098), .A(n1284), 
        .ZN(n1264) );
  AOI221_X1 U661 ( .B1(n1249), .B2(B2[11]), .C1(n1250), .C2(n1085), .A(n1289), 
        .ZN(n1287) );
  NAND2_X1 U849 ( .A1(reg3_reg[1]), .A2(n3704), .ZN(n983) );
  NAND2_X1 U846 ( .A1(reg3_reg[0]), .A2(reg3_reg[1]), .ZN(n988) );
  AOI22_X1 U659 ( .A1(B2[13]), .A2(n985), .B1(n986), .B2(n981), .ZN(n1288) );
  OAI21_X1 U658 ( .B1(B2[12]), .B2(n983), .A(n1288), .ZN(n1275) );
  XNOR2_X1 U657 ( .A(n1287), .B(n1275), .ZN(n1277) );
  XNOR2_X1 U643 ( .A(n1224), .B(n1225), .ZN(n1266) );
  XNOR2_X1 U632 ( .A(n1262), .B(n1233), .ZN(n1032) );
  NOR2_X1 U606 ( .A1(n1233), .A2(n1032), .ZN(n1028) );
  XNOR2_X1 U477 ( .A(n1028), .B(n1029), .ZN(n1026) );
  XNOR2_X1 U652 ( .A(n1265), .B(n1264), .ZN(n1259) );
  AOI22_X1 U681 ( .A1(B2[3]), .A2(n1098), .B1(n1097), .B2(n3827), .ZN(n1311)
         );
  OAI22_X1 U692 ( .A1(B2[11]), .A2(n983), .B1(B2[12]), .B2(n988), .ZN(n1317)
         );
  AOI21_X1 U691 ( .B1(B2[12]), .B2(n985), .A(n1317), .ZN(n1281) );
  AOI22_X1 U651 ( .A1(B2[0]), .A2(n977), .B1(n975), .B2(n989), .ZN(n1278) );
  XNOR2_X1 U666 ( .A(n1260), .B(n1257), .ZN(n1279) );
  AOI222_X1 U631 ( .A1(n1032), .A2(n1033), .B1(n1032), .B2(n1030), .C1(n1033), 
        .C2(n1030), .ZN(p8_C[44]) );
  XNOR2_X1 U649 ( .A(n1258), .B(n1256), .ZN(n1034) );
  AOI22_X1 U695 ( .A1(B2[1]), .A2(n1081), .B1(n1080), .B2(n987), .ZN(n1321) );
  OAI22_X1 U717 ( .A1(B2[11]), .A2(n988), .B1(B2[10]), .B2(n983), .ZN(n1341)
         );
  AOI21_X1 U716 ( .B1(B2[11]), .B2(n985), .A(n1341), .ZN(n1319) );
  XNOR2_X1 U479 ( .A(n1034), .B(n1035), .ZN(p8_S[43]) );
  XNOR2_X1 U715 ( .A(n1318), .B(n1319), .ZN(n1339) );
  XNOR2_X1 U712 ( .A(n1339), .B(n1320), .ZN(n1303) );
  AOI22_X1 U704 ( .A1(B2[4]), .A2(n1123), .B1(n1122), .B2(n1176), .ZN(n1331)
         );
  AOI221_X1 U733 ( .B1(n1148), .B2(B2[4]), .C1(n1149), .C2(n1176), .A(n1349), 
        .ZN(n1333) );
  OAI22_X1 U708 ( .A1(B2[9]), .A2(n983), .B1(B2[7]), .B2(n1212), .ZN(n1337) );
  AOI22_X1 U706 ( .A1(n1333), .A2(n1334), .B1(n1335), .B2(n1336), .ZN(n1332)
         );
  XNOR2_X1 U705 ( .A(n1303), .B(n1332), .ZN(n1305) );
  AOI221_X1 U700 ( .B1(n1107), .B2(B2[3]), .C1(n1108), .C2(n3827), .A(n1330), 
        .ZN(n1300) );
  AOI22_X1 U698 ( .A1(B2[0]), .A2(n1081), .B1(n1080), .B2(n989), .ZN(n1328) );
  XNOR2_X1 U702 ( .A(n1305), .B(n1304), .ZN(n1329) );
  XNOR2_X1 U699 ( .A(n1329), .B(n1300), .ZN(n1302) );
  AOI22_X1 U838 ( .A1(B2[0]), .A2(n1213), .B1(n1212), .B2(n989), .ZN(n1416) );
  AOI221_X1 U837 ( .B1(n1249), .B2(B2[1]), .C1(n1250), .C2(n987), .A(n1416), 
        .ZN(n1076) );
  AOI22_X1 U835 ( .A1(B2[3]), .A2(n985), .B1(n986), .B2(n3827), .ZN(n1415) );
  OAI21_X1 U834 ( .B1(B2[2]), .B2(n983), .A(n1415), .ZN(n1414) );
  AOI221_X1 U850 ( .B1(n1249), .B2(B2[0]), .C1(n1250), .C2(n989), .A(n1421), 
        .ZN(n1078) );
  OAI21_X1 U842 ( .B1(B2[1]), .B2(n983), .A(n1418), .ZN(n1417) );
  NOR2_X1 U840 ( .A1(n1078), .A2(n1079), .ZN(p8_C[32]) );
  OAI221_X1 U823 ( .B1(B2[1]), .B2(n1212), .C1(n987), .C2(n1213), .A(n1411), 
        .ZN(n1071) );
  AOI22_X1 U821 ( .A1(B2[4]), .A2(n985), .B1(n986), .B2(n1176), .ZN(n1410) );
  OAI21_X1 U820 ( .B1(B2[3]), .B2(n983), .A(n1410), .ZN(n1070) );
  XNOR2_X1 U819 ( .A(n1071), .B(n1070), .ZN(n1073) );
  XNOR2_X1 U488 ( .A(n1072), .B(n1073), .ZN(p8_S[34]) );
  NOR2_X1 U832 ( .A1(n1076), .A2(n1077), .ZN(p8_C[33]) );
  AOI22_X1 U811 ( .A1(B2[1]), .A2(n1182), .B1(n1183), .B2(n987), .ZN(n1407) );
  OAI221_X1 U810 ( .B1(B2[0]), .B2(n1168), .C1(n989), .C2(n1169), .A(n1407), 
        .ZN(n1066) );
  AOI221_X1 U816 ( .B1(n1249), .B2(B2[3]), .C1(n1250), .C2(n3827), .A(n1409), 
        .ZN(n1399) );
  OAI21_X1 U812 ( .B1(B2[4]), .B2(n983), .A(n1408), .ZN(n1064) );
  NAND2_X1 U487 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
  NAND2_X1 U807 ( .A1(n1405), .A2(n1406), .ZN(p8_C[35]) );
  NAND2_X1 U485 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
  AOI221_X1 U800 ( .B1(n989), .B2(n1149), .C1(B2[0]), .C2(n1148), .A(n1403), 
        .ZN(n1393) );
  OAI221_X1 U798 ( .B1(B2[1]), .B2(n1168), .C1(n987), .C2(n1169), .A(n1402), 
        .ZN(n1387) );
  OAI22_X1 U782 ( .A1(B2[5]), .A2(n983), .B1(B2[3]), .B2(n1212), .ZN(n1392) );
  AOI221_X1 U781 ( .B1(n985), .B2(B2[6]), .C1(n986), .C2(n1142), .A(n1392), 
        .ZN(n1390) );
  AOI22_X1 U780 ( .A1(B2[4]), .A2(n1249), .B1(n1250), .B2(n1176), .ZN(n1391)
         );
  OAI211_X1 U779 ( .C1(n1213), .C2(n3827), .A(n1390), .B(n1391), .ZN(n1389) );
  OAI21_X1 U778 ( .B1(n1387), .B2(n1388), .A(n1389), .ZN(n1056) );
  AOI22_X1 U794 ( .A1(B2[0]), .A2(n1123), .B1(n1122), .B2(n989), .ZN(n1398) );
  AOI221_X1 U793 ( .B1(n1148), .B2(B2[1]), .C1(n1149), .C2(n987), .A(n1398), 
        .ZN(n1058) );
  AOI22_X1 U792 ( .A1(B2[4]), .A2(n1213), .B1(n1212), .B2(n1176), .ZN(n1397)
         );
  OAI22_X1 U790 ( .A1(B2[6]), .A2(n983), .B1(B2[7]), .B2(n988), .ZN(n1396) );
  AOI21_X1 U789 ( .B1(n985), .B2(B2[7]), .A(n1396), .ZN(n1376) );
  XNOR2_X1 U788 ( .A(n1375), .B(n1376), .ZN(n1394) );
  AOI221_X1 U786 ( .B1(n1182), .B2(B2[3]), .C1(n1183), .C2(n3827), .A(n1395), 
        .ZN(n1377) );
  XNOR2_X1 U785 ( .A(n1394), .B(n1377), .ZN(n1059) );
  OAI21_X1 U797 ( .B1(reg3_reg[7]), .B2(n1063), .A(n1064), .ZN(n1400) );
  OAI22_X1 U795 ( .A1(n1399), .A2(n1400), .B1(n1401), .B2(n3696), .ZN(p8_C[36]) );
  AOI222_X1 U777 ( .A1(n1058), .A2(n1059), .B1(n1058), .B2(n1056), .C1(n1059), 
        .C2(n1056), .ZN(p8_C[37]) );
  AOI22_X1 U776 ( .A1(B2[3]), .A2(n1169), .B1(n1168), .B2(n3827), .ZN(n1386)
         );
  AOI221_X1 U775 ( .B1(n1182), .B2(B2[4]), .C1(n1183), .C2(n1176), .A(n1386), 
        .ZN(n1383) );
  OAI21_X1 U770 ( .B1(B2[7]), .B2(n983), .A(n1384), .ZN(n1370) );
  XNOR2_X1 U769 ( .A(n1371), .B(n1370), .ZN(n1363) );
  XNOR2_X1 U768 ( .A(n1383), .B(n1363), .ZN(n1364) );
  AOI22_X1 U767 ( .A1(B2[1]), .A2(n1123), .B1(n1122), .B2(n987), .ZN(n1382) );
  XNOR2_X1 U758 ( .A(n1362), .B(n1359), .ZN(n1379) );
  AOI222_X1 U755 ( .A1(n1375), .A2(n1376), .B1(n1375), .B2(n1377), .C1(n1376), 
        .C2(n1377), .ZN(n1374) );
  AOI221_X1 U751 ( .B1(n1148), .B2(B2[3]), .C1(n1149), .C2(n3827), .A(n1373), 
        .ZN(n1353) );
  AOI22_X1 U750 ( .A1(B2[4]), .A2(n1169), .B1(n1168), .B2(n1176), .ZN(n1372)
         );
  NAND2_X1 U748 ( .A1(n1370), .A2(n1371), .ZN(n1367) );
  OAI21_X1 U742 ( .B1(B2[8]), .B2(n983), .A(n1368), .ZN(n1350) );
  AOI22_X1 U740 ( .A1(B2[0]), .A2(n1098), .B1(n1097), .B2(n989), .ZN(n1365) );
  NOR2_X1 U753 ( .A1(n1055), .A2(n1054), .ZN(p8_C[38]) );
  AOI22_X1 U737 ( .A1(B2[1]), .A2(n1098), .B1(n1097), .B2(n987), .ZN(n1352) );
  XNOR2_X1 U478 ( .A(n1030), .B(n1031), .ZN(p8_S[44]) );
  AOI222_X1 U648 ( .A1(n1036), .A2(n1037), .B1(n1036), .B2(n1034), .C1(n1037), 
        .C2(n1034), .ZN(p8_C[43]) );
  XNOR2_X1 U476 ( .A(n1022), .B(n1023), .ZN(p8_S[46]) );
  AOI222_X1 U603 ( .A1(n1029), .A2(n1028), .B1(n1029), .B2(n1027), .C1(n1028), 
        .C2(n1027), .ZN(p8_C[45]) );
  XNOR2_X1 U474 ( .A(n1014), .B(n1015), .ZN(p8_S[48]) );
  AOI222_X1 U564 ( .A1(n1020), .A2(n1021), .B1(n1020), .B2(n1018), .C1(n1021), 
        .C2(n1018), .ZN(p8_C[47]) );
  XNOR2_X1 U472 ( .A(n1006), .B(n1007), .ZN(p8_S[50]) );
  AOI222_X1 U532 ( .A1(n1012), .A2(n1013), .B1(n1012), .B2(n1010), .C1(n1013), 
        .C2(n1010), .ZN(p8_C[49]) );
  AOI222_X1 U500 ( .A1(n1093), .A2(n1094), .B1(n1093), .B2(n999), .C1(n1094), 
        .C2(n999), .ZN(p8_C[52]) );
  AOI221_X1 U498 ( .B1(n979), .B2(B2[11]), .C1(n980), .C2(n1085), .A(n1091), 
        .ZN(n995) );
  AOI22_X1 U495 ( .A1(n1086), .A2(n1087), .B1(reg3_reg[13]), .B2(n1088), .ZN(
        n997) );
  XNOR2_X1 U469 ( .A(n994), .B(n997), .ZN(n996) );
  XNOR2_X1 U468 ( .A(n995), .B(n996), .ZN(p8_S[53]) );
  XNOR2_X1 U467 ( .A(n991), .B(n992), .ZN(p8_S[54]) );
  AOI222_X1 U494 ( .A1(n995), .A2(n1083), .B1(n995), .B2(n997), .C1(n1083), 
        .C2(n997), .ZN(p8_C[53]) );
  AOI22_X1 U462 ( .A1(B2[13]), .A2(n979), .B1(n980), .B2(n981), .ZN(n978) );
  OAI221_X1 U461 ( .B1(B2[12]), .B2(n975), .C1(n976), .C2(n977), .A(n978), 
        .ZN(p8_final_product2_26_) );
  NOR2_X1 U1475 ( .A1(n3674), .A2(n3724), .ZN(n1881) );
  OAI21_X1 U1473 ( .B1(reg1_reg[11]), .B2(reg1_reg[12]), .A(n1876), .ZN(n2208)
         );
  AOI221_X1 U1293 ( .B1(n1878), .B2(B0[11]), .C1(n1879), .C2(n1984), .A(n1990), 
        .ZN(n1894) );
  OAI21_X1 U1524 ( .B1(reg1_reg[9]), .B2(reg1_reg[10]), .A(n1980), .ZN(n2246)
         );
  AOI22_X1 U1292 ( .A1(B0[13]), .A2(n1988), .B1(n1989), .B2(n1880), .ZN(n1981)
         );
  OAI221_X1 U1291 ( .B1(B0[12]), .B2(n1979), .C1(n1875), .C2(n1980), .A(n1981), 
        .ZN(n1982) );
  OAI21_X1 U1560 ( .B1(reg1_reg[7]), .B2(reg1_reg[8]), .A(n1997), .ZN(n2281)
         );
  AOI22_X1 U1308 ( .A1(B0[13]), .A2(n2006), .B1(n2007), .B2(n1880), .ZN(n1998)
         );
  OAI221_X1 U1297 ( .B1(B0[13]), .B2(n1996), .C1(n1880), .C2(n1997), .A(n1998), 
        .ZN(n1995) );
  AOI22_X1 U1299 ( .A1(B0[12]), .A2(n1988), .B1(n1989), .B2(n1875), .ZN(n1999)
         );
  OAI221_X1 U1298 ( .B1(B0[11]), .B2(n1979), .C1(n1984), .C2(n1980), .A(n1999), 
        .ZN(n1986) );
  AOI22_X1 U1290 ( .A1(n1985), .A2(n1986), .B1(reg1_reg[13]), .B2(n1987), .ZN(
        n1896) );
  XNOR2_X1 U1264 ( .A(n1893), .B(n1896), .ZN(n1895) );
  OAI221_X1 U1307 ( .B1(B0[12]), .B2(n1996), .C1(n1875), .C2(n1997), .A(n1998), 
        .ZN(n1899) );
  AOI221_X1 U1309 ( .B1(n1988), .B2(B0[11]), .C1(n1989), .C2(n1984), .A(n2008), 
        .ZN(n2002) );
  AOI22_X1 U1305 ( .A1(B0[8]), .A2(n1876), .B1(n1874), .B2(n2005), .ZN(n2004)
         );
  OAI22_X1 U1301 ( .A1(n2000), .A2(n2001), .B1(n2002), .B2(n1899), .ZN(n1900)
         );
  OAI21_X1 U1601 ( .B1(reg1_reg[6]), .B2(reg1_reg[5]), .A(n2022), .ZN(n2304)
         );
  AOI22_X1 U1357 ( .A1(B0[11]), .A2(n2022), .B1(n2021), .B2(n1984), .ZN(n2070)
         );
  AOI221_X1 U1356 ( .B1(n2047), .B2(B0[12]), .C1(n2048), .C2(n1875), .A(n2070), 
        .ZN(n2049) );
  OAI21_X1 U1626 ( .B1(reg1_reg[3]), .B2(reg1_reg[4]), .A(n2068), .ZN(n2313)
         );
  AOI22_X1 U1371 ( .A1(B0[13]), .A2(n2081), .B1(n2082), .B2(n1880), .ZN(n2069)
         );
  OAI221_X1 U1355 ( .B1(B0[13]), .B2(n2067), .C1(n1880), .C2(n2068), .A(n2069), 
        .ZN(n2050) );
  XNOR2_X1 U1354 ( .A(n2049), .B(n2050), .ZN(n2051) );
  OAI22_X1 U1339 ( .A1(n2049), .A2(n2050), .B1(n2051), .B2(n2052), .ZN(n2031)
         );
  AOI22_X1 U1338 ( .A1(B0[13]), .A2(n2047), .B1(n2048), .B2(n1880), .ZN(n2023)
         );
  OAI221_X1 U1337 ( .B1(B0[12]), .B2(n2021), .C1(n1875), .C2(n2022), .A(n2023), 
        .ZN(n2011) );
  AOI221_X1 U1335 ( .B1(n2006), .B2(B0[11]), .C1(n2007), .C2(n1984), .A(n2046), 
        .ZN(n2033) );
  AOI22_X1 U1334 ( .A1(B0[8]), .A2(n1980), .B1(n1979), .B2(n2005), .ZN(n2045)
         );
  XNOR2_X1 U1351 ( .A(n2051), .B(n2052), .ZN(n2038) );
  AOI221_X1 U1348 ( .B1(n1988), .B2(B0[8]), .C1(n1989), .C2(n2005), .A(n2064), 
        .ZN(n2039) );
  AOI221_X1 U1372 ( .B1(n2047), .B2(B0[11]), .C1(n2048), .C2(n1984), .A(n2083), 
        .ZN(n2071) );
  OAI221_X1 U1370 ( .B1(B0[12]), .B2(n2067), .C1(n1875), .C2(n2068), .A(n2069), 
        .ZN(n2035) );
  XNOR2_X1 U1369 ( .A(n2071), .B(n2035), .ZN(n2072) );
  OAI221_X1 U1367 ( .B1(B0[8]), .B2(n1996), .C1(n2005), .C2(n1997), .A(n2080), 
        .ZN(n2079) );
  OAI22_X1 U1358 ( .A1(n2071), .A2(n2035), .B1(n2072), .B2(n2073), .ZN(n2065)
         );
  XNOR2_X1 U1350 ( .A(n2065), .B(n2038), .ZN(n2040) );
  XNOR2_X1 U1347 ( .A(n2040), .B(n2039), .ZN(n2060) );
  AOI22_X1 U1328 ( .A1(n2034), .A2(n2035), .B1(n2036), .B2(n2037), .ZN(n1909)
         );
  AOI222_X1 U1327 ( .A1(n1911), .A2(n1912), .B1(n1911), .B2(n1909), .C1(n1912), 
        .C2(n1909), .ZN(p6_C[49]) );
  AOI22_X1 U1322 ( .A1(B0[11]), .A2(n1997), .B1(n1996), .B2(n1984), .ZN(n2024)
         );
  AOI221_X1 U1321 ( .B1(n2006), .B2(B0[12]), .C1(n2007), .C2(n1875), .A(n2024), 
        .ZN(n2020) );
  OAI221_X1 U1320 ( .B1(B0[13]), .B2(n2021), .C1(n1880), .C2(n2022), .A(n2023), 
        .ZN(n2014) );
  XNOR2_X1 U1319 ( .A(n2020), .B(n2014), .ZN(n2015) );
  XNOR2_X1 U1316 ( .A(n2015), .B(n2013), .ZN(n2016) );
  AOI22_X1 U1315 ( .A1(B0[8]), .A2(n1878), .B1(n1879), .B2(n2005), .ZN(n2018)
         );
  AOI22_X1 U1324 ( .A1(n2029), .A2(n2030), .B1(n2031), .B2(n2032), .ZN(n1907)
         );
  AOI22_X1 U1323 ( .A1(n2025), .A2(n2026), .B1(n2027), .B2(n2028), .ZN(n1908)
         );
  XNOR2_X1 U1267 ( .A(n1905), .B(n1906), .ZN(p6_S[50]) );
  XNOR2_X1 U1268 ( .A(n1909), .B(n1910), .ZN(p6_S[49]) );
  OAI21_X1 U1652 ( .B1(reg1_reg[1]), .B2(reg1_reg[2]), .A(n2112), .ZN(n2322)
         );
  NAND2_X1 U1648 ( .A1(reg1_reg[3]), .A2(n2322), .ZN(n2111) );
  AOI22_X1 U1421 ( .A1(B0[13]), .A2(n2148), .B1(n2149), .B2(n1880), .ZN(n2113)
         );
  OAI221_X1 U1391 ( .B1(B0[13]), .B2(n2111), .C1(n1880), .C2(n2112), .A(n2113), 
        .ZN(n2087) );
  AOI22_X1 U1390 ( .A1(B0[12]), .A2(n2081), .B1(n2082), .B2(n1875), .ZN(n2110)
         );
  OAI221_X1 U1389 ( .B1(B0[11]), .B2(n2067), .C1(n1984), .C2(n2068), .A(n2110), 
        .ZN(n2109) );
  NAND2_X1 U1375 ( .A1(n2084), .A2(n2087), .ZN(n2086) );
  OAI21_X1 U1374 ( .B1(n2084), .B2(n2085), .A(n2086), .ZN(n2078) );
  AOI221_X1 U1392 ( .B1(n2006), .B2(B0[8]), .C1(n2007), .C2(n2005), .A(n2114), 
        .ZN(n2089) );
  AOI22_X1 U1376 ( .A1(n2088), .A2(n2089), .B1(n2090), .B2(n2091), .ZN(n2057)
         );
  AOI22_X1 U1341 ( .A1(n2056), .A2(n2057), .B1(n2058), .B2(n2059), .ZN(n1916)
         );
  AOI22_X1 U1362 ( .A1(B0[4]), .A2(n1876), .B1(n1874), .B2(n2075), .ZN(n2074)
         );
  XNOR2_X1 U1363 ( .A(n2076), .B(n2054), .ZN(n2055) );
  AOI222_X1 U1340 ( .A1(n1915), .A2(n1916), .B1(n1915), .B2(n1913), .C1(n1916), 
        .C2(n1913), .ZN(p6_C[48]) );
  XNOR2_X1 U1360 ( .A(n2055), .B(n2053), .ZN(n1917) );
  AOI22_X1 U1415 ( .A1(B0[8]), .A2(n2022), .B1(n2021), .B2(n2005), .ZN(n2145)
         );
  OAI221_X1 U1420 ( .B1(B0[12]), .B2(n2111), .C1(n1875), .C2(n2112), .A(n2113), 
        .ZN(n2095) );
  AOI221_X1 U1422 ( .B1(n2081), .B2(B0[11]), .C1(n2082), .C2(n1984), .A(n2150), 
        .ZN(n2147) );
  XNOR2_X1 U1419 ( .A(n2147), .B(n2095), .ZN(n2105) );
  AOI22_X1 U1412 ( .A1(B0[4]), .A2(n1980), .B1(n1979), .B2(n2075), .ZN(n2143)
         );
  XNOR2_X1 U1416 ( .A(n2105), .B(n2118), .ZN(n2144) );
  XNOR2_X1 U1413 ( .A(n2144), .B(n2104), .ZN(n2119) );
  AOI22_X1 U1380 ( .A1(n2097), .A2(n2098), .B1(n2099), .B2(n2100), .ZN(n1919)
         );
  AOI22_X1 U1395 ( .A1(B0[4]), .A2(n1878), .B1(n1879), .B2(n2075), .ZN(n2116)
         );
  OAI221_X1 U1394 ( .B1(B0[3]), .B2(n1874), .C1(n2115), .C2(n1876), .A(n2116), 
        .ZN(n2094) );
  AOI22_X1 U1379 ( .A1(n2093), .A2(n2094), .B1(n2095), .B2(n2096), .ZN(n1920)
         );
  XNOR2_X1 U1270 ( .A(n1917), .B(n1918), .ZN(p6_S[47]) );
  XNOR2_X1 U1410 ( .A(n2119), .B(n2117), .ZN(n2125) );
  NAND2_X1 U1644 ( .A1(n3715), .A2(reg1_reg[0]), .ZN(n1889) );
  AOI22_X1 U1435 ( .A1(B0[13]), .A2(n1884), .B1(reg1_reg[1]), .B2(n1880), .ZN(
        n2151) );
  AOI22_X1 U1433 ( .A1(B0[11]), .A2(n2112), .B1(n2111), .B2(n1984), .ZN(n2170)
         );
  AOI221_X1 U1432 ( .B1(n2148), .B2(B0[12]), .C1(n2149), .C2(n1875), .A(n2170), 
        .ZN(n2169) );
  OAI22_X1 U1424 ( .A1(n2151), .A2(n2152), .B1(n2153), .B2(n2154), .ZN(n2142)
         );
  AOI22_X1 U1442 ( .A1(B0[3]), .A2(n1980), .B1(n1979), .B2(n2115), .ZN(n2173)
         );
  AOI22_X1 U1440 ( .A1(B0[1]), .A2(n1876), .B1(n1874), .B2(n1886), .ZN(n2172)
         );
  NOR2_X1 U1409 ( .A1(n2123), .A2(n2124), .ZN(n2141) );
  XNOR2_X1 U1408 ( .A(n2127), .B(n2141), .ZN(n2135) );
  XNOR2_X1 U1404 ( .A(n2135), .B(n2126), .ZN(n2120) );
  AOI22_X1 U1403 ( .A1(B0[3]), .A2(n1878), .B1(n1879), .B2(n2115), .ZN(n2134)
         );
  OAI21_X1 U1397 ( .B1(n2123), .B2(n2124), .A(n2120), .ZN(n2122) );
  OAI21_X1 U1396 ( .B1(n2120), .B2(n2121), .A(n2122), .ZN(n1924) );
  AOI222_X1 U1383 ( .A1(n1923), .A2(n1924), .B1(n1923), .B2(n1921), .C1(n1924), 
        .C2(n1921), .ZN(p6_C[46]) );
  OAI221_X1 U1448 ( .B1(B0[4]), .B2(n1996), .C1(n2075), .C2(n1997), .A(n2183), 
        .ZN(n2163) );
  AOI221_X1 U1456 ( .B1(n2148), .B2(B0[11]), .C1(n2149), .C2(n1984), .A(n2188), 
        .ZN(n2186) );
  NAND2_X1 U1645 ( .A1(reg1_reg[1]), .A2(n3722), .ZN(n1882) );
  NAND2_X1 U1642 ( .A1(reg1_reg[0]), .A2(reg1_reg[1]), .ZN(n1887) );
  AOI22_X1 U1454 ( .A1(B0[13]), .A2(n1884), .B1(n1885), .B2(n1880), .ZN(n2187)
         );
  OAI21_X1 U1453 ( .B1(B0[12]), .B2(n1882), .A(n2187), .ZN(n2174) );
  XNOR2_X1 U1452 ( .A(n2186), .B(n2174), .ZN(n2176) );
  OAI221_X1 U1450 ( .B1(B0[8]), .B2(n2067), .C1(n2005), .C2(n2068), .A(n2185), 
        .ZN(n2175) );
  XNOR2_X1 U1427 ( .A(n2161), .B(n2132), .ZN(n1931) );
  XNOR2_X1 U1272 ( .A(n1927), .B(n1928), .ZN(n1925) );
  XNOR2_X1 U1447 ( .A(n2164), .B(n2163), .ZN(n2158) );
  AOI22_X1 U1477 ( .A1(B0[3]), .A2(n1997), .B1(n1996), .B2(n2115), .ZN(n2212)
         );
  OAI22_X1 U1488 ( .A1(B0[11]), .A2(n1882), .B1(B0[12]), .B2(n1887), .ZN(n2218) );
  AOI21_X1 U1487 ( .B1(B0[12]), .B2(n1884), .A(n2218), .ZN(n2180) );
  AOI22_X1 U1446 ( .A1(B0[0]), .A2(n1876), .B1(n1874), .B2(n1888), .ZN(n2177)
         );
  XNOR2_X1 U1461 ( .A(n2159), .B(n2156), .ZN(n2178) );
  XNOR2_X1 U1444 ( .A(n2157), .B(n2155), .ZN(n1933) );
  AOI22_X1 U1491 ( .A1(B0[1]), .A2(n1980), .B1(n1979), .B2(n1886), .ZN(n2222)
         );
  OAI22_X1 U1513 ( .A1(B0[11]), .A2(n1887), .B1(B0[10]), .B2(n1882), .ZN(n2241) );
  AOI21_X1 U1512 ( .B1(B0[11]), .B2(n1884), .A(n2241), .ZN(n2220) );
  XNOR2_X1 U1274 ( .A(n1933), .B(n1934), .ZN(p6_S[43]) );
  XNOR2_X1 U1508 ( .A(n2239), .B(n2221), .ZN(n2202) );
  AOI22_X1 U1500 ( .A1(B0[4]), .A2(n2022), .B1(n2021), .B2(n2075), .ZN(n2231)
         );
  AOI221_X1 U1506 ( .B1(B0[8]), .B2(n2148), .C1(n2149), .C2(n2005), .A(n2238), 
        .ZN(n2235) );
  OAI22_X1 U1504 ( .A1(B0[9]), .A2(n1882), .B1(B0[7]), .B2(n2111), .ZN(n2237)
         );
  AOI22_X1 U1502 ( .A1(n2233), .A2(n2234), .B1(n2235), .B2(n2236), .ZN(n2232)
         );
  XNOR2_X1 U1501 ( .A(n2202), .B(n2232), .ZN(n2204) );
  AOI22_X1 U1494 ( .A1(B0[0]), .A2(n1980), .B1(n1979), .B2(n1888), .ZN(n2228)
         );
  AOI22_X1 U1634 ( .A1(B0[0]), .A2(n2112), .B1(n2111), .B2(n1888), .ZN(n2316)
         );
  AOI221_X1 U1633 ( .B1(n2148), .B2(B0[1]), .C1(n2149), .C2(n1886), .A(n2316), 
        .ZN(n1975) );
  AOI22_X1 U1631 ( .A1(B0[3]), .A2(n1884), .B1(n1885), .B2(n2115), .ZN(n2315)
         );
  OAI21_X1 U1630 ( .B1(B0[2]), .B2(n1882), .A(n2315), .ZN(n2314) );
  NOR2_X1 U1636 ( .A1(n1977), .A2(n1978), .ZN(p6_C[32]) );
  OAI221_X1 U1619 ( .B1(B0[1]), .B2(n2111), .C1(n1886), .C2(n2112), .A(n2311), 
        .ZN(n1970) );
  AOI22_X1 U1617 ( .A1(B0[4]), .A2(n1884), .B1(n1885), .B2(n2075), .ZN(n2310)
         );
  OAI21_X1 U1616 ( .B1(B0[3]), .B2(n1882), .A(n2310), .ZN(n1969) );
  XNOR2_X1 U1615 ( .A(n1970), .B(n1969), .ZN(n1972) );
  XNOR2_X1 U1283 ( .A(n1971), .B(n1972), .ZN(p6_S[34]) );
  NOR2_X1 U1628 ( .A1(n1975), .A2(n1976), .ZN(p6_C[33]) );
  AOI22_X1 U1607 ( .A1(B0[1]), .A2(n2081), .B1(n2082), .B2(n1886), .ZN(n2307)
         );
  OAI221_X1 U1606 ( .B1(B0[0]), .B2(n2067), .C1(n1888), .C2(n2068), .A(n2307), 
        .ZN(n1965) );
  OAI21_X1 U1608 ( .B1(B0[4]), .B2(n1882), .A(n2308), .ZN(n1963) );
  NAND2_X1 U1603 ( .A1(n2305), .A2(n2306), .ZN(p6_C[35]) );
  NAND2_X1 U1280 ( .A1(n1963), .A2(n1964), .ZN(n1961) );
  OAI221_X1 U1594 ( .B1(B0[1]), .B2(n2067), .C1(n1886), .C2(n2068), .A(n2302), 
        .ZN(n2287) );
  OAI22_X1 U1578 ( .A1(B0[5]), .A2(n1882), .B1(B0[3]), .B2(n2111), .ZN(n2292)
         );
  AOI22_X1 U1576 ( .A1(B0[4]), .A2(n2148), .B1(n2149), .B2(n2075), .ZN(n2291)
         );
  OAI211_X1 U1575 ( .C1(n2112), .C2(n2115), .A(n2290), .B(n2291), .ZN(n2289)
         );
  OAI21_X1 U1574 ( .B1(n2287), .B2(n2288), .A(n2289), .ZN(n1955) );
  AOI22_X1 U1590 ( .A1(B0[0]), .A2(n2022), .B1(n2021), .B2(n1888), .ZN(n2298)
         );
  AOI221_X1 U1589 ( .B1(n2047), .B2(B0[1]), .C1(n2048), .C2(n1886), .A(n2298), 
        .ZN(n1957) );
  AOI22_X1 U1588 ( .A1(B0[4]), .A2(n2112), .B1(n2111), .B2(n2075), .ZN(n2297)
         );
  OAI22_X1 U1586 ( .A1(B0[6]), .A2(n1882), .B1(B0[7]), .B2(n1887), .ZN(n2296)
         );
  AOI21_X1 U1585 ( .B1(n1884), .B2(B0[7]), .A(n2296), .ZN(n2276) );
  XNOR2_X1 U1584 ( .A(n2275), .B(n2276), .ZN(n2294) );
  AOI221_X1 U1582 ( .B1(n2081), .B2(B0[3]), .C1(n2082), .C2(n2115), .A(n2295), 
        .ZN(n2277) );
  XNOR2_X1 U1581 ( .A(n2294), .B(n2277), .ZN(n1958) );
  OAI21_X1 U1593 ( .B1(reg1_reg[7]), .B2(n1962), .A(n1963), .ZN(n2300) );
  OAI22_X1 U1591 ( .A1(n2299), .A2(n2300), .B1(n2301), .B2(n3710), .ZN(
        p6_C[36]) );
  AOI222_X1 U1573 ( .A1(n1957), .A2(n1958), .B1(n1957), .B2(n1955), .C1(n1958), 
        .C2(n1955), .ZN(p6_C[37]) );
  AOI222_X1 U1551 ( .A1(n2275), .A2(n2276), .B1(n2275), .B2(n2277), .C1(n2276), 
        .C2(n2277), .ZN(n2274) );
  AOI22_X1 U1572 ( .A1(B0[3]), .A2(n2068), .B1(n2067), .B2(n2115), .ZN(n2286)
         );
  AOI221_X1 U1571 ( .B1(n2081), .B2(B0[4]), .C1(n2082), .C2(n2075), .A(n2286), 
        .ZN(n2283) );
  XNOR2_X1 U1564 ( .A(n2283), .B(n2263), .ZN(n2264) );
  AOI22_X1 U1563 ( .A1(B0[1]), .A2(n2022), .B1(n2021), .B2(n1886), .ZN(n2282)
         );
  AOI22_X1 U1552 ( .A1(reg1_reg[9]), .A2(n2278), .B1(n2261), .B2(n3713), .ZN(
        n1954) );
  AOI22_X1 U1546 ( .A1(B0[4]), .A2(n2068), .B1(n2067), .B2(n2075), .ZN(n2272)
         );
  AOI22_X1 U1536 ( .A1(B0[0]), .A2(n1997), .B1(n1996), .B2(n1888), .ZN(n2265)
         );
  NOR2_X1 U1549 ( .A1(n1954), .A2(n1953), .ZN(p6_C[38]) );
  AOI22_X1 U1533 ( .A1(B0[1]), .A2(n1997), .B1(n1996), .B2(n1886), .ZN(n2252)
         );
  AOI222_X1 U1443 ( .A1(n1935), .A2(n1936), .B1(n1935), .B2(n1933), .C1(n1936), 
        .C2(n1933), .ZN(p6_C[43]) );
  XNOR2_X1 U1271 ( .A(n1921), .B(n1922), .ZN(p6_S[46]) );
  AOI222_X1 U1398 ( .A1(n1928), .A2(n1927), .B1(n1928), .B2(n1926), .C1(n1927), 
        .C2(n1926), .ZN(p6_C[45]) );
  XNOR2_X1 U1269 ( .A(n1913), .B(n1914), .ZN(p6_S[48]) );
  AOI222_X1 U1359 ( .A1(n1919), .A2(n1920), .B1(n1919), .B2(n1917), .C1(n1920), 
        .C2(n1917), .ZN(p6_C[47]) );
  AOI222_X1 U1313 ( .A1(n1907), .A2(n1908), .B1(n1907), .B2(n1905), .C1(n1908), 
        .C2(n1905), .ZN(p6_C[50]) );
  XNOR2_X1 U1303 ( .A(n2000), .B(n2001), .ZN(n1901) );
  AOI22_X1 U1311 ( .A1(n2009), .A2(n2010), .B1(n2011), .B2(n2012), .ZN(n1904)
         );
  XNOR2_X1 U1266 ( .A(n1901), .B(n1902), .ZN(p6_S[51]) );
  XNOR2_X1 U1265 ( .A(n1897), .B(n1898), .ZN(p6_S[52]) );
  AOI222_X1 U1302 ( .A1(n1903), .A2(n1904), .B1(n1903), .B2(n1901), .C1(n1904), 
        .C2(n1901), .ZN(p6_C[51]) );
  AOI22_X1 U1288 ( .A1(B0[11]), .A2(n1876), .B1(n1874), .B2(n1984), .ZN(n1983)
         );
  AOI221_X1 U1287 ( .B1(n1878), .B2(B0[12]), .C1(n1879), .C2(n1875), .A(n1983), 
        .ZN(n1892) );
  OAI221_X1 U1285 ( .B1(B0[13]), .B2(n1979), .C1(n1880), .C2(n1980), .A(n1981), 
        .ZN(n1891) );
  XNOR2_X1 U1262 ( .A(n1890), .B(n1891), .ZN(p6_S[54]) );
  AOI222_X1 U1289 ( .A1(n1894), .A2(n1982), .B1(n1894), .B2(n1896), .C1(n1982), 
        .C2(n1896), .ZN(p6_C[53]) );
  AOI22_X1 U1258 ( .A1(B0[13]), .A2(n1878), .B1(n1879), .B2(n1880), .ZN(n1877)
         );
  OAI221_X1 U1257 ( .B1(B0[12]), .B2(n1874), .C1(n1875), .C2(n1876), .A(n1877), 
        .ZN(p6_final_product2_26_) );
  NOR2_X1 U50 ( .A1(n1881), .A2(n1878), .ZN(n513) );
  AOI22_X1 U2089 ( .A1(reg4[10]), .A2(n2776), .B1(n2774), .B2(n3682), .ZN(
        n2890) );
  AOI221_X1 U2088 ( .B1(n2778), .B2(reg4[11]), .C1(n2779), .C2(n3671), .A(
        n2890), .ZN(n2794) );
  AOI22_X1 U2087 ( .A1(reg4[13]), .A2(n2888), .B1(n2889), .B2(n3676), .ZN(
        n2881) );
  OAI221_X1 U2086 ( .B1(reg4[12]), .B2(n2879), .C1(n3679), .C2(n2880), .A(
        n2881), .ZN(n2882) );
  AOI22_X1 U2103 ( .A1(reg4[13]), .A2(n2906), .B1(n2907), .B2(n3676), .ZN(
        n2898) );
  AOI22_X1 U2094 ( .A1(reg4[12]), .A2(n2888), .B1(n2889), .B2(n3679), .ZN(
        n2899) );
  OAI221_X1 U2093 ( .B1(reg4[11]), .B2(n2879), .C1(n3671), .C2(n2880), .A(
        n2899), .ZN(n2886) );
  AOI22_X1 U2085 ( .A1(n2885), .A2(n2886), .B1(A2[13]), .B2(n2887), .ZN(n2796)
         );
  XNOR2_X1 U2058 ( .A(n2793), .B(n2796), .ZN(n2795) );
  XNOR2_X1 U2057 ( .A(n2794), .B(n2795), .ZN(p10_S[53]) );
  AOI22_X1 U2105 ( .A1(reg4[10]), .A2(n2880), .B1(n2879), .B2(n3682), .ZN(
        n2908) );
  AOI221_X1 U2104 ( .B1(n2888), .B2(reg4[11]), .C1(n2889), .C2(n3671), .A(
        n2908), .ZN(n2902) );
  AOI22_X1 U2100 ( .A1(reg4[8]), .A2(n2776), .B1(n2774), .B2(n3667), .ZN(n2904) );
  AOI221_X1 U2099 ( .B1(n2778), .B2(reg4[9]), .C1(n2779), .C2(n3681), .A(n2904), .ZN(n2901) );
  OAI22_X1 U2096 ( .A1(n2900), .A2(n2901), .B1(n2902), .B2(n2799), .ZN(n2800)
         );
  AOI22_X1 U2166 ( .A1(reg4[13]), .A2(n2984), .B1(n2985), .B2(n3676), .ZN(
        n2969) );
  XNOR2_X1 U2149 ( .A(n2949), .B(n2950), .ZN(n2951) );
  AOI221_X1 U2147 ( .B1(n2906), .B2(reg4[10]), .C1(n2907), .C2(n3682), .A(
        n2966), .ZN(n2952) );
  OAI22_X1 U2134 ( .A1(n2949), .A2(n2950), .B1(n2951), .B2(n2952), .ZN(n2931)
         );
  AOI22_X1 U2133 ( .A1(reg4[13]), .A2(n2947), .B1(n2948), .B2(n3676), .ZN(
        n2923) );
  AOI221_X1 U2130 ( .B1(n2906), .B2(reg4[11]), .C1(n2907), .C2(n3671), .A(
        n2946), .ZN(n2933) );
  AOI22_X1 U2129 ( .A1(reg4[8]), .A2(n2880), .B1(n2879), .B2(n3667), .ZN(n2945) );
  AOI221_X1 U2128 ( .B1(n2888), .B2(reg4[9]), .C1(n2889), .C2(n3681), .A(n2945), .ZN(n2944) );
  AOI22_X1 U2125 ( .A1(reg4[7]), .A2(n2778), .B1(n2779), .B2(n3672), .ZN(n2942) );
  OAI221_X1 U2124 ( .B1(reg4[6]), .B2(n2774), .C1(n3678), .C2(n2776), .A(n2942), .ZN(n2926) );
  XNOR2_X1 U2146 ( .A(n2951), .B(n2952), .ZN(n2938) );
  AOI22_X1 U2144 ( .A1(reg4[7]), .A2(n2880), .B1(n2879), .B2(n3672), .ZN(n2964) );
  AOI221_X1 U2143 ( .B1(n2888), .B2(reg4[8]), .C1(n2889), .C2(n3667), .A(n2964), .ZN(n2939) );
  XNOR2_X1 U2164 ( .A(n2971), .B(n2935), .ZN(n2972) );
  AOI22_X1 U2163 ( .A1(reg4[9]), .A2(n2906), .B1(n2907), .B2(n3681), .ZN(n2983) );
  OAI22_X1 U2153 ( .A1(n2971), .A2(n2935), .B1(n2972), .B2(n2973), .ZN(n2965)
         );
  XNOR2_X1 U2145 ( .A(n2965), .B(n2938), .ZN(n2940) );
  XNOR2_X1 U2142 ( .A(n2940), .B(n2939), .ZN(n2960) );
  AOI22_X1 U2141 ( .A1(reg4[5]), .A2(n2776), .B1(n2774), .B2(n3664), .ZN(n2962) );
  AOI22_X1 U2123 ( .A1(n2934), .A2(n2935), .B1(n2936), .B2(n2937), .ZN(n2809)
         );
  AOI222_X1 U2122 ( .A1(n2811), .A2(n2812), .B1(n2811), .B2(n2809), .C1(n2812), 
        .C2(n2809), .ZN(p10_C[49]) );
  AOI221_X1 U2116 ( .B1(n2906), .B2(reg4[12]), .C1(n2907), .C2(n3679), .A(
        n2924), .ZN(n2920) );
  XNOR2_X1 U2114 ( .A(n2920), .B(n2914), .ZN(n2915) );
  AOI22_X1 U2113 ( .A1(reg4[9]), .A2(n2880), .B1(n2879), .B2(n3681), .ZN(n2919) );
  AOI221_X1 U2112 ( .B1(n2888), .B2(reg4[10]), .C1(n2889), .C2(n3682), .A(
        n2919), .ZN(n2913) );
  XNOR2_X1 U2111 ( .A(n2915), .B(n2913), .ZN(n2916) );
  AOI22_X1 U2110 ( .A1(reg4[8]), .A2(n2778), .B1(n2779), .B2(n3667), .ZN(n2918) );
  OAI221_X1 U2109 ( .B1(reg4[7]), .B2(n2774), .C1(n3672), .C2(n2776), .A(n2918), .ZN(n2910) );
  AOI22_X1 U2119 ( .A1(n2929), .A2(n2930), .B1(n2931), .B2(n2932), .ZN(n2807)
         );
  AOI22_X1 U2118 ( .A1(n2925), .A2(n2926), .B1(n2927), .B2(n2928), .ZN(n2808)
         );
  XNOR2_X1 U2061 ( .A(n2805), .B(n2806), .ZN(p10_S[50]) );
  XNOR2_X1 U2062 ( .A(n2809), .B(n2810), .ZN(p10_S[49]) );
  AOI22_X1 U2210 ( .A1(reg4[13]), .A2(n3047), .B1(n3048), .B2(n3676), .ZN(
        n3010) );
  AOI221_X1 U2182 ( .B1(n2984), .B2(reg4[12]), .C1(n2985), .C2(n3679), .A(
        n3011), .ZN(n3007) );
  XNOR2_X1 U2180 ( .A(n3007), .B(n2980), .ZN(n2981) );
  AOI221_X1 U2185 ( .B1(n2906), .B2(reg4[8]), .C1(n2907), .C2(n3667), .A(n3012), .ZN(n2988) );
  XNOR2_X1 U2184 ( .A(n2979), .B(n2988), .ZN(n3006) );
  AOI22_X1 U2179 ( .A1(reg4[6]), .A2(n2888), .B1(n2889), .B2(n3678), .ZN(n3005) );
  OAI221_X1 U2178 ( .B1(reg4[5]), .B2(n2879), .C1(n3664), .C2(n2880), .A(n3005), .ZN(n2991) );
  AOI22_X1 U2169 ( .A1(n2987), .A2(n2988), .B1(n2989), .B2(n2990), .ZN(n2957)
         );
  AOI22_X1 U2136 ( .A1(n2956), .A2(n2957), .B1(n2958), .B2(n2959), .ZN(n2816)
         );
  AOI22_X1 U2157 ( .A1(reg4[4]), .A2(n2776), .B1(n2774), .B2(n3668), .ZN(n2974) );
  AOI221_X1 U2156 ( .B1(n2778), .B2(reg4[5]), .C1(n2779), .C2(n3664), .A(n2974), .ZN(n2953) );
  AOI22_X1 U2160 ( .A1(reg4[6]), .A2(n2880), .B1(n2879), .B2(n3678), .ZN(n2977) );
  AOI221_X1 U2159 ( .B1(n2888), .B2(reg4[7]), .C1(n2889), .C2(n3672), .A(n2977), .ZN(n2954) );
  XNOR2_X1 U2158 ( .A(n2976), .B(n2954), .ZN(n2955) );
  AOI221_X1 U2211 ( .B1(n2984), .B2(reg4[11]), .C1(n2985), .C2(n3671), .A(
        n3049), .ZN(n3046) );
  XNOR2_X1 U2208 ( .A(n3046), .B(n2994), .ZN(n3004) );
  AOI22_X1 U2206 ( .A1(reg4[4]), .A2(n2880), .B1(n2879), .B2(n3668), .ZN(n3044) );
  AOI221_X1 U2214 ( .B1(n2906), .B2(reg4[7]), .C1(n2907), .C2(n3672), .A(n3050), .ZN(n3017) );
  XNOR2_X1 U2213 ( .A(n3003), .B(n3017), .ZN(n3045) );
  XNOR2_X1 U2207 ( .A(n3045), .B(n3004), .ZN(n3018) );
  AOI22_X1 U2173 ( .A1(n2996), .A2(n2997), .B1(n2998), .B2(n2999), .ZN(n2819)
         );
  AOI22_X1 U2190 ( .A1(reg4[4]), .A2(n2778), .B1(n2779), .B2(n3668), .ZN(n3015) );
  OAI221_X1 U2189 ( .B1(reg4[3]), .B2(n2774), .C1(n3665), .C2(n2776), .A(n3015), .ZN(n2993) );
  AOI22_X1 U2172 ( .A1(n2992), .A2(n2993), .B1(n2994), .B2(n2995), .ZN(n2820)
         );
  XNOR2_X1 U2155 ( .A(n2955), .B(n2953), .ZN(n2817) );
  AOI222_X1 U2154 ( .A1(n2819), .A2(n2820), .B1(n2819), .B2(n2817), .C1(n2820), 
        .C2(n2817), .ZN(p10_C[47]) );
  XNOR2_X1 U2063 ( .A(n2813), .B(n2814), .ZN(p10_S[48]) );
  XNOR2_X1 U2064 ( .A(n2817), .B(n2818), .ZN(p10_S[47]) );
  XNOR2_X1 U2204 ( .A(n3018), .B(n3016), .ZN(n3024) );
  AOI221_X1 U2229 ( .B1(n2947), .B2(reg4[8]), .C1(n2948), .C2(n3667), .A(n3070), .ZN(n3069) );
  AOI22_X1 U2227 ( .A1(reg4[13]), .A2(n2784), .B1(A2[1]), .B2(n3676), .ZN(
        n3068) );
  AOI22_X1 U2225 ( .A1(reg4[12]), .A2(n3047), .B1(n3048), .B2(n3679), .ZN(
        n3067) );
  AOI221_X1 U2222 ( .B1(n2984), .B2(reg4[10]), .C1(n2985), .C2(n3682), .A(
        n3065), .ZN(n3041) );
  AOI22_X1 U2221 ( .A1(reg4[6]), .A2(n2906), .B1(n2907), .B2(n3678), .ZN(n3063) );
  AOI22_X1 U2200 ( .A1(n3035), .A2(n3036), .B1(n3037), .B2(n3038), .ZN(n3025)
         );
  AOI22_X1 U2235 ( .A1(reg4[3]), .A2(n2880), .B1(n2879), .B2(n3665), .ZN(n3072) );
  AOI22_X1 U2233 ( .A1(reg4[1]), .A2(n2776), .B1(n2774), .B2(n3666), .ZN(n3071) );
  NOR2_X1 U2203 ( .A1(n3022), .A2(n3023), .ZN(n3039) );
  XNOR2_X1 U2202 ( .A(n3026), .B(n3039), .ZN(n3034) );
  XNOR2_X1 U2199 ( .A(n3034), .B(n3025), .ZN(n3019) );
  AOI22_X1 U2198 ( .A1(reg4[3]), .A2(n2778), .B1(n2779), .B2(n3665), .ZN(n3033) );
  OAI221_X1 U2197 ( .B1(reg4[2]), .B2(n2774), .C1(n3673), .C2(n2776), .A(n3033), .ZN(n3020) );
  OAI21_X1 U2192 ( .B1(n3022), .B2(n3023), .A(n3019), .ZN(n3021) );
  OAI21_X1 U2191 ( .B1(n3019), .B2(n3020), .A(n3021), .ZN(n2824) );
  AOI221_X1 U2323 ( .B1(n2906), .B2(reg4[2]), .C1(n2907), .C2(n3673), .A(n3150), .ZN(n3124) );
  NAND2_X1 U2428 ( .A1(A2[0]), .A2(A2[1]), .ZN(n2787) );
  AOI22_X1 U2330 ( .A1(reg4[9]), .A2(n2784), .B1(n2785), .B2(n3681), .ZN(n3166) );
  OAI21_X1 U2329 ( .B1(reg4[8]), .B2(n2782), .A(n3166), .ZN(n3148) );
  AOI221_X1 U2320 ( .B1(n2947), .B2(reg4[4]), .C1(n2948), .C2(n3668), .A(n3147), .ZN(n3131) );
  AOI221_X1 U2318 ( .B1(n2984), .B2(reg4[6]), .C1(n2985), .C2(n3678), .A(n3146), .ZN(n3132) );
  AOI221_X1 U2304 ( .B1(n3047), .B2(reg4[9]), .C1(n3048), .C2(n3681), .A(n3140), .ZN(n3116) );
  OAI22_X1 U2303 ( .A1(reg4[11]), .A2(n2787), .B1(reg4[10]), .B2(n2782), .ZN(
        n3139) );
  AOI21_X1 U2302 ( .B1(reg4[11]), .B2(n2784), .A(n3139), .ZN(n3117) );
  XNOR2_X1 U2301 ( .A(n3116), .B(n3117), .ZN(n3137) );
  AOI221_X1 U2299 ( .B1(n2984), .B2(reg4[7]), .C1(n2985), .C2(n3672), .A(n3138), .ZN(n3118) );
  XNOR2_X1 U2298 ( .A(n3137), .B(n3118), .ZN(n3101) );
  NOR2_X1 U2297 ( .A1(n3009), .A2(n3672), .ZN(n3136) );
  AOI221_X1 U2296 ( .B1(reg4[8]), .B2(n3047), .C1(n3048), .C2(n3667), .A(n3136), .ZN(n3133) );
  AOI221_X1 U2294 ( .B1(n2785), .B2(n3682), .C1(n2784), .C2(reg4[10]), .A(
        n3135), .ZN(n3134) );
  XNOR2_X1 U2292 ( .A(n3101), .B(n3130), .ZN(n3103) );
  XNOR2_X1 U2289 ( .A(n3103), .B(n3102), .ZN(n3127) );
  AOI221_X1 U2287 ( .B1(n2906), .B2(reg4[3]), .C1(n2907), .C2(n3665), .A(n3128), .ZN(n3098) );
  XNOR2_X1 U2286 ( .A(n3127), .B(n3098), .ZN(n3100) );
  AOI22_X1 U2285 ( .A1(reg4[0]), .A2(n2880), .B1(n2879), .B2(n3670), .ZN(n3126) );
  XNOR2_X1 U2070 ( .A(n2841), .B(n2842), .ZN(p10_S[41]) );
  AOI221_X1 U2334 ( .B1(n2984), .B2(reg4[5]), .C1(n2985), .C2(n3664), .A(n3170), .ZN(n3155) );
  AOI22_X1 U2357 ( .A1(reg4[8]), .A2(n2784), .B1(n2785), .B2(n3667), .ZN(n3182) );
  OAI21_X1 U2356 ( .B1(reg4[7]), .B2(n2782), .A(n3182), .ZN(n3168) );
  AOI22_X1 U2359 ( .A1(reg4[6]), .A2(n3047), .B1(n3048), .B2(n3678), .ZN(n3183) );
  NAND2_X1 U2333 ( .A1(n3168), .A2(n3169), .ZN(n3165) );
  AOI221_X1 U2336 ( .B1(n2947), .B2(reg4[3]), .C1(n2948), .C2(n3665), .A(n3171), .ZN(n3151) );
  AOI221_X1 U2326 ( .B1(n2906), .B2(reg4[1]), .C1(n2907), .C2(n3666), .A(n3163), .ZN(n3152) );
  AOI221_X1 U2344 ( .B1(n2906), .B2(reg4[0]), .C1(n2907), .C2(n3670), .A(n3178), .ZN(n3157) );
  AOI221_X1 U2360 ( .B1(n2984), .B2(reg4[4]), .C1(n2985), .C2(n3668), .A(n3184), .ZN(n3181) );
  XNOR2_X1 U2355 ( .A(n3169), .B(n3168), .ZN(n3161) );
  XNOR2_X1 U2354 ( .A(n3181), .B(n3161), .ZN(n3162) );
  AOI221_X1 U2352 ( .B1(n2947), .B2(reg4[2]), .C1(n2948), .C2(n3673), .A(n3180), .ZN(n3160) );
  XNOR2_X1 U2343 ( .A(n3160), .B(n3157), .ZN(n3177) );
  AOI221_X1 U2377 ( .B1(n3047), .B2(reg4[5]), .C1(n3048), .C2(n3664), .A(n3197), .ZN(n3173) );
  OAI22_X1 U2376 ( .A1(reg4[6]), .A2(n2782), .B1(reg4[7]), .B2(n2787), .ZN(
        n3196) );
  AOI21_X1 U2375 ( .B1(n2784), .B2(reg4[7]), .A(n3196), .ZN(n3174) );
  AOI221_X1 U2372 ( .B1(n2984), .B2(reg4[3]), .C1(n2985), .C2(n3665), .A(n3195), .ZN(n3175) );
  AOI222_X1 U2340 ( .A1(n3173), .A2(n3174), .B1(n3173), .B2(n3175), .C1(n3174), 
        .C2(n3175), .ZN(n3172) );
  AOI22_X1 U2368 ( .A1(n3664), .A2(n3192), .B1(n3665), .B2(n3709), .ZN(n3191)
         );
  OAI221_X1 U2367 ( .B1(n2789), .B2(n3678), .C1(n2787), .C2(reg4[6]), .A(n3191), .ZN(n3190) );
  AOI221_X1 U2366 ( .B1(n3668), .B2(n3048), .C1(reg4[4]), .C2(n3047), .A(n3190), .ZN(n3186) );
  AOI221_X1 U2385 ( .B1(n2984), .B2(reg4[2]), .C1(n2985), .C2(n3673), .A(n3201), .ZN(n3189) );
  AOI221_X1 U2364 ( .B1(n3186), .B2(n3665), .C1(n3186), .C2(n3009), .A(n3187), 
        .ZN(n2855) );
  XNOR2_X1 U2374 ( .A(n3173), .B(n3174), .ZN(n3194) );
  XNOR2_X1 U2371 ( .A(n3194), .B(n3175), .ZN(n2858) );
  AOI22_X1 U2402 ( .A1(reg4[5]), .A2(n2784), .B1(n2785), .B2(n3664), .ZN(n3207) );
  OAI21_X1 U2401 ( .B1(reg4[4]), .B2(n2782), .A(n3207), .ZN(n2863) );
  NAND2_X1 U2382 ( .A1(A2[7]), .A2(n2861), .ZN(n3200) );
  NAND2_X1 U2381 ( .A1(n3199), .A2(n3200), .ZN(p10_C[36]) );
  AOI22_X1 U2399 ( .A1(reg4[1]), .A2(n2984), .B1(n2985), .B2(n3666), .ZN(n3206) );
  AOI22_X1 U2410 ( .A1(reg4[4]), .A2(n2784), .B1(n2785), .B2(n3668), .ZN(n3210) );
  OAI21_X1 U2409 ( .B1(reg4[3]), .B2(n2782), .A(n3210), .ZN(n2870) );
  NAND2_X1 U2077 ( .A1(n2869), .A2(n2870), .ZN(n2868) );
  AOI221_X1 U2422 ( .B1(n3047), .B2(reg4[1]), .C1(n3048), .C2(n3666), .A(n3216), .ZN(n2875) );
  AOI22_X1 U2420 ( .A1(reg4[3]), .A2(n2784), .B1(n2785), .B2(n3665), .ZN(n3215) );
  OAI21_X1 U2419 ( .B1(reg4[2]), .B2(n2782), .A(n3215), .ZN(n3214) );
  AOI221_X1 U2432 ( .B1(n3670), .B2(n3048), .C1(reg4[0]), .C2(n3047), .A(n3709), .ZN(n2878) );
  OAI22_X1 U2427 ( .A1(reg4[1]), .A2(n2782), .B1(reg4[2]), .B2(n2787), .ZN(
        n3217) );
  AOI21_X1 U2426 ( .B1(n2784), .B2(reg4[2]), .A(n3217), .ZN(n2877) );
  OAI221_X1 U2055 ( .B1(reg4[0]), .B2(n2787), .C1(n3670), .C2(n2789), .A(n2782), .ZN(\p10/final_product1[0] ) );
  NOR2_X1 U2417 ( .A1(n2875), .A2(n2876), .ZN(p10_C[33]) );
  NAND2_X1 U2395 ( .A1(n3204), .A2(n3205), .ZN(p10_C[35]) );
  AOI222_X1 U2362 ( .A1(n2857), .A2(n2858), .B1(n2857), .B2(n3185), .C1(n2858), 
        .C2(n3185), .ZN(p10_C[37]) );
  AOI222_X1 U2283 ( .A1(n2843), .A2(n2844), .B1(n2843), .B2(n2841), .C1(n2844), 
        .C2(n2841), .ZN(p10_C[41]) );
  OAI22_X1 U2277 ( .A1(reg4[11]), .A2(n2782), .B1(reg4[12]), .B2(n2787), .ZN(
        n3114) );
  AOI21_X1 U2276 ( .B1(reg4[12]), .B2(n2784), .A(n3114), .ZN(n3080) );
  AOI221_X1 U2270 ( .B1(n2984), .B2(reg4[8]), .C1(n2985), .C2(n3667), .A(n3111), .ZN(n3081) );
  AOI221_X1 U2267 ( .B1(n2906), .B2(reg4[4]), .C1(n2907), .C2(n3668), .A(n3109), .ZN(n3091) );
  AOI22_X1 U2282 ( .A1(reg4[1]), .A2(n2880), .B1(n2879), .B2(n3666), .ZN(n3119) );
  AOI22_X1 U2254 ( .A1(reg4[7]), .A2(n2947), .B1(n2948), .B2(n3672), .ZN(n3089) );
  AOI221_X1 U2251 ( .B1(n3047), .B2(reg4[11]), .C1(n3048), .C2(n3671), .A(
        n3088), .ZN(n3086) );
  AOI22_X1 U2250 ( .A1(reg4[13]), .A2(n2784), .B1(n2785), .B2(n3676), .ZN(
        n3087) );
  OAI21_X1 U2249 ( .B1(reg4[12]), .B2(n2782), .A(n3087), .ZN(n3073) );
  XNOR2_X1 U2248 ( .A(n3086), .B(n3073), .ZN(n3075) );
  AOI22_X1 U2247 ( .A1(reg4[9]), .A2(n2984), .B1(n2985), .B2(n3681), .ZN(n3085) );
  AOI22_X1 U2245 ( .A1(reg4[5]), .A2(n2906), .B1(n2907), .B2(n3664), .ZN(n3083) );
  XNOR2_X1 U2243 ( .A(n3061), .B(n3060), .ZN(n3055) );
  XNOR2_X1 U2242 ( .A(n3056), .B(n3057), .ZN(n3077) );
  AOI22_X1 U2241 ( .A1(reg4[2]), .A2(n2880), .B1(n2879), .B2(n3673), .ZN(n3078) );
  AOI22_X1 U2239 ( .A1(reg4[0]), .A2(n2776), .B1(n2774), .B2(n3670), .ZN(n3076) );
  XNOR2_X1 U2237 ( .A(n3054), .B(n3052), .ZN(n2833) );
  XNOR2_X1 U2068 ( .A(n2833), .B(n2834), .ZN(p10_S[43]) );
  XNOR2_X1 U2231 ( .A(n3022), .B(n3023), .ZN(n3062) );
  XNOR2_X1 U2219 ( .A(n3058), .B(n3031), .ZN(n2831) );
  AOI222_X1 U2236 ( .A1(n2835), .A2(n2836), .B1(n2835), .B2(n2833), .C1(n2836), 
        .C2(n2833), .ZN(p10_C[43]) );
  XNOR2_X1 U2066 ( .A(n2827), .B(n2828), .ZN(n2825) );
  AOI22_X1 U2194 ( .A1(n3027), .A2(n3028), .B1(n3029), .B2(n3030), .ZN(n2826)
         );
  AOI222_X1 U2218 ( .A1(n2831), .A2(n2832), .B1(n2831), .B2(n2829), .C1(n2832), 
        .C2(n2829), .ZN(p10_C[44]) );
  XNOR2_X1 U2065 ( .A(n2821), .B(n2822), .ZN(p10_S[46]) );
  AOI222_X1 U2193 ( .A1(n2828), .A2(n2827), .B1(n2828), .B2(n2826), .C1(n2827), 
        .C2(n2826), .ZN(p10_C[45]) );
  XNOR2_X1 U2098 ( .A(n2900), .B(n2901), .ZN(n2801) );
  AOI22_X1 U2106 ( .A1(n2909), .A2(n2910), .B1(n2911), .B2(n2912), .ZN(n2804)
         );
  XNOR2_X1 U2060 ( .A(n2801), .B(n2802), .ZN(p10_S[51]) );
  AOI222_X1 U2108 ( .A1(n2807), .A2(n2808), .B1(n2807), .B2(n2805), .C1(n2808), 
        .C2(n2805), .ZN(p10_C[50]) );
  XNOR2_X1 U2059 ( .A(n2797), .B(n2798), .ZN(p10_S[52]) );
  AOI222_X1 U2097 ( .A1(n2803), .A2(n2804), .B1(n2803), .B2(n2801), .C1(n2804), 
        .C2(n2801), .ZN(p10_C[51]) );
  AOI22_X1 U2083 ( .A1(reg4[11]), .A2(n2776), .B1(n2774), .B2(n3671), .ZN(
        n2883) );
  AOI221_X1 U2082 ( .B1(n2778), .B2(reg4[12]), .C1(n2779), .C2(n3679), .A(
        n2883), .ZN(n2792) );
  OAI221_X1 U2080 ( .B1(reg4[13]), .B2(n2879), .C1(n3676), .C2(n2880), .A(
        n2881), .ZN(n2791) );
  AOI222_X1 U2079 ( .A1(n2792), .A2(n2793), .B1(n2792), .B2(n2791), .C1(n2793), 
        .C2(n2791), .ZN(p10_C[54]) );
  AOI22_X1 U2051 ( .A1(reg4[13]), .A2(n2778), .B1(n2779), .B2(n3676), .ZN(
        n2777) );
  OAI221_X1 U2050 ( .B1(reg4[12]), .B2(n2774), .C1(n3679), .C2(n2776), .A(
        n2777), .ZN(p10_final_product2_26_) );
  NOR2_X1 U58 ( .A1(n2781), .A2(n2778), .ZN(n521) );
  NAND2_X1 U2469 ( .A1(n3230), .A2(n3728), .ZN(n3229) );
  NAND2_X1 U2466 ( .A1(n3225), .A2(n3729), .ZN(n3224) );
  NAND2_X1 U2463 ( .A1(n3222), .A2(n3730), .ZN(n3244) );
  NOR2_X1 U2459 ( .A1(reg7[10]), .A2(n3244), .ZN(n3242) );
  NAND2_X1 U2458 ( .A1(n3242), .A2(n3748), .ZN(n3241) );
  NOR2_X1 U2457 ( .A1(n3241), .A2(reg7[12]), .ZN(n3240) );
  NOR2_X1 U2462 ( .A1(reg7[10]), .A2(reg7[9]), .ZN(n3245) );
  AOI22_X1 U2461 ( .A1(n3244), .A2(reg7[10]), .B1(n3222), .B2(n3245), .ZN(
        SUB1_N10) );
  AOI22_X1 U2440 ( .A1(reg7[9]), .A2(n3221), .B1(n3222), .B2(n3730), .ZN(
        SUB1_N9) );
  NOR2_X1 U2443 ( .A1(reg7[8]), .A2(reg7[7]), .ZN(n3226) );
  AOI22_X1 U2442 ( .A1(n3224), .A2(reg7[8]), .B1(n3225), .B2(n3226), .ZN(
        SUB1_N8) );
  AOI22_X1 U2444 ( .A1(n3225), .A2(n3729), .B1(reg7[7]), .B2(n3228), .ZN(
        SUB1_N7) );
  NOR2_X1 U2447 ( .A1(reg7[6]), .A2(reg7[5]), .ZN(n3231) );
  AOI22_X1 U2446 ( .A1(n3229), .A2(reg7[6]), .B1(n3230), .B2(n3231), .ZN(
        SUB1_N6) );
  AOI22_X1 U2448 ( .A1(n3230), .A2(n3728), .B1(reg7[5]), .B2(n3233), .ZN(
        SUB1_N5) );
  NOR2_X1 U2451 ( .A1(reg7[4]), .A2(reg7[3]), .ZN(n3236) );
  AOI22_X1 U2450 ( .A1(n3234), .A2(reg7[4]), .B1(n3235), .B2(n3236), .ZN(
        SUB1_N4) );
  AOI22_X1 U2452 ( .A1(n3235), .A2(n3727), .B1(reg7[3]), .B2(n3238), .ZN(
        SUB1_N3) );
  NOR2_X1 U2455 ( .A1(reg7[1]), .A2(reg7[0]), .ZN(n3239) );
  XNOR2_X1 U2454 ( .A(n3239), .B(reg7[2]), .ZN(SUB1_N2) );
  AOI22_X1 U2475 ( .A1(reg7[0]), .A2(reg7[1]), .B1(n3731), .B2(n3707), .ZN(
        SUB1_N1) );
  NAND2_X1 U2757 ( .A1(VIN), .A2(w[13]), .ZN(n3327) );
  OAI21_X1 U2756 ( .B1(VIN), .B2(n3680), .A(n3327), .ZN(REG11_n48) );
  OAI21_X1 U2616 ( .B1(VIN), .B2(n3757), .A(n3327), .ZN(REGISTER1_n48) );
  NAND2_X1 U2505 ( .A1(VIN), .A2(ff[13]), .ZN(n3261) );
  OAI21_X1 U2504 ( .B1(VIN), .B2(REGISTER_out_n75), .A(n3261), .ZN(
        REGISTER_out_n48) );
  NAND2_X1 U2754 ( .A1(VIN), .A2(w[12]), .ZN(n3326) );
  OAI21_X1 U2753 ( .B1(VIN), .B2(n3690), .A(n3326), .ZN(REG11_n49) );
  OAI21_X1 U2614 ( .B1(VIN), .B2(n3724), .A(n3326), .ZN(REGISTER1_n49) );
  NAND2_X1 U2503 ( .A1(VIN), .A2(ff[12]), .ZN(n3260) );
  OAI21_X1 U2502 ( .B1(VIN), .B2(REGISTER_out_n74), .A(n3260), .ZN(
        REGISTER_out_n49) );
  NAND2_X1 U2751 ( .A1(VIN), .A2(w[11]), .ZN(n3325) );
  OAI21_X1 U2750 ( .B1(VIN), .B2(n3686), .A(n3325), .ZN(REG11_n50) );
  OAI21_X1 U2612 ( .B1(VIN), .B2(n3674), .A(n3325), .ZN(REGISTER1_n50) );
  NAND2_X1 U2501 ( .A1(VIN), .A2(ff[11]), .ZN(n3259) );
  OAI21_X1 U2500 ( .B1(VIN), .B2(REGISTER_out_n73), .A(n3259), .ZN(
        REGISTER_out_n50) );
  NAND2_X1 U2748 ( .A1(VIN), .A2(w[10]), .ZN(n3324) );
  OAI21_X1 U2747 ( .B1(VIN), .B2(n3693), .A(n3324), .ZN(REG11_n51) );
  OAI21_X1 U2610 ( .B1(VIN), .B2(n3749), .A(n3324), .ZN(REGISTER1_n51) );
  NAND2_X1 U2499 ( .A1(VIN), .A2(ff[10]), .ZN(n3258) );
  OAI21_X1 U2498 ( .B1(VIN), .B2(REGISTER_out_n72), .A(n3258), .ZN(
        REGISTER_out_n51) );
  NAND2_X1 U2745 ( .A1(VIN), .A2(w[9]), .ZN(n3322) );
  OAI21_X1 U2744 ( .B1(VIN), .B2(n3691), .A(n3322), .ZN(REG11_n52) );
  OAI21_X1 U2608 ( .B1(VIN), .B2(n3713), .A(n3322), .ZN(REGISTER1_n52) );
  NAND2_X1 U2497 ( .A1(VIN), .A2(ff[9]), .ZN(n3257) );
  OAI21_X1 U2496 ( .B1(VIN), .B2(REGISTER_out_n71), .A(n3257), .ZN(
        REGISTER_out_n52) );
  NAND2_X1 U2742 ( .A1(VIN), .A2(w[8]), .ZN(n3321) );
  OAI21_X1 U2741 ( .B1(VIN), .B2(n3683), .A(n3321), .ZN(REG11_n53) );
  OAI21_X1 U2606 ( .B1(VIN), .B2(n3750), .A(n3321), .ZN(REGISTER1_n53) );
  NAND2_X1 U2495 ( .A1(VIN), .A2(ff[8]), .ZN(n3256) );
  OAI21_X1 U2494 ( .B1(VIN), .B2(REGISTER_out_n70), .A(n3256), .ZN(
        REGISTER_out_n53) );
  NAND2_X1 U2739 ( .A1(VIN), .A2(w[7]), .ZN(n3319) );
  OAI21_X1 U2738 ( .B1(VIN), .B2(n3688), .A(n3319), .ZN(REG11_n54) );
  OAI21_X1 U2604 ( .B1(VIN), .B2(n3710), .A(n3319), .ZN(REGISTER1_n54) );
  NAND2_X1 U2493 ( .A1(VIN), .A2(ff[7]), .ZN(n3255) );
  OAI21_X1 U2492 ( .B1(VIN), .B2(REGISTER_out_n69), .A(n3255), .ZN(
        REGISTER_out_n54) );
  NAND2_X1 U2736 ( .A1(VIN), .A2(w[6]), .ZN(n3318) );
  OAI21_X1 U2735 ( .B1(VIN), .B2(n3687), .A(n3318), .ZN(REG11_n55) );
  OAI21_X1 U2602 ( .B1(VIN), .B2(n3759), .A(n3318), .ZN(REGISTER1_n55) );
  NAND2_X1 U2491 ( .A1(VIN), .A2(ff[6]), .ZN(n3254) );
  OAI21_X1 U2490 ( .B1(VIN), .B2(REGISTER_out_n68), .A(n3254), .ZN(
        REGISTER_out_n55) );
  NAND2_X1 U2733 ( .A1(VIN), .A2(w[5]), .ZN(n3316) );
  OAI21_X1 U2732 ( .B1(VIN), .B2(n3677), .A(n3316), .ZN(REG11_n56) );
  OAI21_X1 U2600 ( .B1(VIN), .B2(n3711), .A(n3316), .ZN(REGISTER1_n56) );
  NAND2_X1 U2489 ( .A1(VIN), .A2(ff[5]), .ZN(n3253) );
  OAI21_X1 U2488 ( .B1(VIN), .B2(REGISTER_out_n67), .A(n3253), .ZN(
        REGISTER_out_n56) );
  NAND2_X1 U2730 ( .A1(VIN), .A2(w[4]), .ZN(n3315) );
  OAI21_X1 U2729 ( .B1(VIN), .B2(n3685), .A(n3315), .ZN(REG11_n57) );
  OAI21_X1 U2598 ( .B1(VIN), .B2(n3751), .A(n3315), .ZN(REGISTER1_n57) );
  NAND2_X1 U2487 ( .A1(VIN), .A2(ff[4]), .ZN(n3252) );
  OAI21_X1 U2486 ( .B1(VIN), .B2(REGISTER_out_n66), .A(n3252), .ZN(
        REGISTER_out_n57) );
  NAND2_X1 U2727 ( .A1(VIN), .A2(w[3]), .ZN(n3313) );
  OAI21_X1 U2726 ( .B1(VIN), .B2(n3669), .A(n3313), .ZN(REG11_n58) );
  OAI21_X1 U2596 ( .B1(VIN), .B2(n3717), .A(n3313), .ZN(REGISTER1_n58) );
  NAND2_X1 U2485 ( .A1(VIN), .A2(ff[3]), .ZN(n3251) );
  OAI21_X1 U2484 ( .B1(VIN), .B2(REGISTER_out_n65), .A(n3251), .ZN(
        REGISTER_out_n58) );
  OAI21_X1 U2652 ( .B1(VIN), .B2(n3665), .A(n3294), .ZN(REG31_n58) );
  OAI21_X1 U2656 ( .B1(VIN), .B2(n3664), .A(n3297), .ZN(REG31_n56) );
  OAI21_X1 U2672 ( .B1(VIN), .B2(n3676), .A(n3308), .ZN(REG31_n48) );
  OAI21_X1 U2654 ( .B1(VIN), .B2(n3668), .A(n3296), .ZN(REG31_n57) );
  OAI21_X1 U2648 ( .B1(VIN), .B2(n3666), .A(n3291), .ZN(REG31_n60) );
  OAI21_X1 U2646 ( .B1(VIN), .B2(n3670), .A(n3290), .ZN(REG31_n61) );
  OAI21_X1 U2658 ( .B1(VIN), .B2(n3678), .A(n3299), .ZN(REG31_n55) );
  OAI21_X1 U2660 ( .B1(VIN), .B2(n3672), .A(n3300), .ZN(REG31_n54) );
  OAI21_X1 U2664 ( .B1(VIN), .B2(n3681), .A(n3303), .ZN(REG31_n52) );
  OAI21_X1 U2662 ( .B1(VIN), .B2(n3667), .A(n3302), .ZN(REG31_n53) );
  OAI21_X1 U2650 ( .B1(VIN), .B2(n3673), .A(n3293), .ZN(REG31_n59) );
  OAI21_X1 U2666 ( .B1(VIN), .B2(n3682), .A(n3305), .ZN(REG31_n51) );
  OAI21_X1 U2668 ( .B1(VIN), .B2(n3671), .A(n3306), .ZN(REG31_n50) );
  OAI21_X1 U2670 ( .B1(VIN), .B2(n3679), .A(n3307), .ZN(REG31_n49) );
  NAND2_X1 U2724 ( .A1(VIN), .A2(w[2]), .ZN(n3312) );
  OAI21_X1 U2723 ( .B1(VIN), .B2(n3692), .A(n3312), .ZN(REG11_n59) );
  OAI21_X1 U2594 ( .B1(VIN), .B2(n3752), .A(n3312), .ZN(REGISTER1_n59) );
  OAI21_X1 U2588 ( .B1(VIN), .B2(n3758), .A(n3308), .ZN(REGISTER2_n48) );
  OAI21_X1 U2572 ( .B1(VIN), .B2(n3712), .A(n3297), .ZN(REGISTER2_n56) );
  OAI21_X1 U2576 ( .B1(VIN), .B2(n3714), .A(n3300), .ZN(REGISTER2_n54) );
  OAI21_X1 U2580 ( .B1(VIN), .B2(n3719), .A(n3303), .ZN(REGISTER2_n52) );
  OAI21_X1 U2695 ( .B1(VIN), .B2(n3734), .A(n3300), .ZN(REG21_n54) );
  OAI21_X1 U2677 ( .B1(VIN), .B2(n3737), .A(n3291), .ZN(REG21_n60) );
  OAI21_X1 U2564 ( .B1(VIN), .B2(n3716), .A(n3291), .ZN(REGISTER2_n60) );
  OAI21_X1 U2683 ( .B1(VIN), .B2(n3736), .A(n3294), .ZN(REG21_n58) );
  OAI21_X1 U2701 ( .B1(VIN), .B2(n3733), .A(n3303), .ZN(REG21_n52) );
  OAI21_X1 U2689 ( .B1(VIN), .B2(n3735), .A(n3297), .ZN(REG21_n56) );
  OAI21_X1 U2713 ( .B1(VIN), .B2(n3708), .A(n3308), .ZN(REG21_n48) );
  OAI21_X1 U2674 ( .B1(VIN), .B2(n3738), .A(n3290), .ZN(REG21_n61) );
  OAI21_X1 U2562 ( .B1(VIN), .B2(n3723), .A(n3290), .ZN(REGISTER2_n61) );
  OAI21_X1 U2584 ( .B1(VIN), .B2(n3694), .A(n3306), .ZN(REGISTER2_n50) );
  OAI21_X1 U2568 ( .B1(VIN), .B2(n3718), .A(n3294), .ZN(REGISTER2_n58) );
  OAI21_X1 U2570 ( .B1(VIN), .B2(n3755), .A(n3296), .ZN(REGISTER2_n57) );
  OAI21_X1 U2686 ( .B1(VIN), .B2(n3766), .A(n3296), .ZN(REG21_n57) );
  OAI21_X1 U2566 ( .B1(VIN), .B2(n3756), .A(n3293), .ZN(REGISTER2_n59) );
  OAI21_X1 U2680 ( .B1(VIN), .B2(n3767), .A(n3293), .ZN(REG21_n59) );
  OAI21_X1 U2574 ( .B1(VIN), .B2(n3760), .A(n3299), .ZN(REGISTER2_n55) );
  OAI21_X1 U2692 ( .B1(VIN), .B2(n3765), .A(n3299), .ZN(REG21_n55) );
  OAI21_X1 U2704 ( .B1(VIN), .B2(n3763), .A(n3305), .ZN(REG21_n51) );
  OAI21_X1 U2582 ( .B1(VIN), .B2(n3753), .A(n3305), .ZN(REGISTER2_n51) );
  OAI21_X1 U2707 ( .B1(VIN), .B2(n3732), .A(n3306), .ZN(REG21_n50) );
  OAI21_X1 U2586 ( .B1(VIN), .B2(n3725), .A(n3307), .ZN(REGISTER2_n49) );
  OAI21_X1 U2710 ( .B1(VIN), .B2(n3762), .A(n3307), .ZN(REG21_n49) );
  OAI21_X1 U2698 ( .B1(VIN), .B2(n3764), .A(n3302), .ZN(REG21_n53) );
  OAI21_X1 U2578 ( .B1(VIN), .B2(n3754), .A(n3302), .ZN(REGISTER2_n53) );
  OAI22_X1 U2523 ( .A1(n3852), .A2(reg5[8]), .B1(reg4_reg[8]), .B2(VIN), .ZN(
        n3270) );
  OAI22_X1 U2515 ( .A1(n3849), .A2(reg5[4]), .B1(reg4_reg[4]), .B2(VIN), .ZN(
        n3266) );
  OAI22_X1 U2547 ( .A1(n3849), .A2(reg3[6]), .B1(reg3_reg[6]), .B2(VIN), .ZN(
        n3282) );
  OAI22_X1 U2519 ( .A1(n3849), .A2(reg5[6]), .B1(reg4_reg[6]), .B2(VIN), .ZN(
        n3268) );
  OAI22_X1 U2559 ( .A1(n3849), .A2(reg3[12]), .B1(reg3_reg[12]), .B2(VIN), 
        .ZN(n3288) );
  OAI22_X1 U2527 ( .A1(n3847), .A2(reg5[10]), .B1(reg4_reg[10]), .B2(VIN), 
        .ZN(n3272) );
  OAI22_X1 U2539 ( .A1(n3847), .A2(reg3[2]), .B1(reg3_reg[2]), .B2(VIN), .ZN(
        n3278) );
  OAI22_X1 U2555 ( .A1(n3846), .A2(reg3[10]), .B1(reg3_reg[10]), .B2(VIN), 
        .ZN(n3286) );
  OAI22_X1 U2543 ( .A1(n3847), .A2(reg3[4]), .B1(reg3_reg[4]), .B2(VIN), .ZN(
        n3280) );
  OAI22_X1 U2511 ( .A1(n3849), .A2(reg5[2]), .B1(reg4_reg[2]), .B2(VIN), .ZN(
        n3264) );
  OAI22_X1 U2551 ( .A1(n3851), .A2(reg3[8]), .B1(reg3_reg[8]), .B2(VIN), .ZN(
        n3284) );
  NAND2_X1 U2721 ( .A1(VIN), .A2(w[1]), .ZN(n3310) );
  OAI21_X1 U2720 ( .B1(VIN), .B2(n3684), .A(n3310), .ZN(REG11_n60) );
  OAI21_X1 U2717 ( .B1(VIN), .B2(n3689), .A(n3309), .ZN(REG11_n61) );
  OAI21_X1 U2590 ( .B1(VIN), .B2(n3722), .A(n3309), .ZN(REGISTER1_n61) );
  OAI21_X1 U2592 ( .B1(VIN), .B2(n3715), .A(n3310), .ZN(REGISTER1_n60) );
  AOI22_X1 U2628 ( .A1(VIN), .A2(n3664), .B1(n3744), .B2(n3851), .ZN(REG41_n56) );
  AOI22_X1 U2624 ( .A1(VIN), .A2(n3665), .B1(n3745), .B2(n3850), .ZN(REG41_n58) );
  AOI22_X1 U2644 ( .A1(VIN), .A2(n3676), .B1(n3739), .B2(n3850), .ZN(REG41_n48) );
  AOI22_X1 U2620 ( .A1(VIN), .A2(n3666), .B1(n3746), .B2(n3850), .ZN(REG41_n60) );
  AOI22_X1 U2626 ( .A1(VIN), .A2(n3668), .B1(n3771), .B2(n3851), .ZN(REG41_n57) );
  AOI22_X1 U2634 ( .A1(VIN), .A2(n3667), .B1(n3769), .B2(n3848), .ZN(REG41_n53) );
  AOI22_X1 U2630 ( .A1(VIN), .A2(n3678), .B1(n3770), .B2(n3847), .ZN(REG41_n55) );
  AOI22_X1 U2618 ( .A1(VIN), .A2(n3670), .B1(n3747), .B2(n3850), .ZN(REG41_n61) );
  AOI22_X1 U2636 ( .A1(VIN), .A2(n3681), .B1(n3742), .B2(n3847), .ZN(REG41_n52) );
  AOI22_X1 U2642 ( .A1(VIN), .A2(n3679), .B1(n3740), .B2(n3846), .ZN(REG41_n49) );
  AOI22_X1 U2640 ( .A1(VIN), .A2(n3671), .B1(n3741), .B2(n3848), .ZN(REG41_n50) );
  AOI22_X1 U2632 ( .A1(VIN), .A2(n3672), .B1(n3743), .B2(n3848), .ZN(REG41_n54) );
  AOI22_X1 U2638 ( .A1(VIN), .A2(n3682), .B1(n3768), .B2(n3846), .ZN(REG41_n51) );
  AOI22_X1 U2622 ( .A1(VIN), .A2(n3673), .B1(n3772), .B2(n3852), .ZN(REG41_n59) );
  AOI22_X1 U2512 ( .A1(VIN), .A2(n3745), .B1(n3703), .B2(n3848), .ZN(
        REGISTER4_n58) );
  AOI22_X1 U2552 ( .A1(VIN), .A2(n3733), .B1(n3721), .B2(n3851), .ZN(
        REGISTER3_n52) );
  AOI22_X1 U2516 ( .A1(VIN), .A2(n3744), .B1(n3699), .B2(n3852), .ZN(
        REGISTER4_n56) );
  AOI22_X1 U2544 ( .A1(VIN), .A2(n3735), .B1(n3698), .B2(n3846), .ZN(
        REGISTER3_n56) );
  AOI22_X1 U2540 ( .A1(VIN), .A2(n3736), .B1(n3702), .B2(n3846), .ZN(
        REGISTER3_n58) );
  AOI22_X1 U2548 ( .A1(VIN), .A2(n3734), .B1(n3696), .B2(n3849), .ZN(
        REGISTER3_n54) );
  AOI22_X1 U2520 ( .A1(VIN), .A2(n3743), .B1(n3697), .B2(n3848), .ZN(
        REGISTER4_n54) );
  AOI22_X1 U2508 ( .A1(VIN), .A2(n3746), .B1(n3701), .B2(n3846), .ZN(
        REGISTER4_n60) );
  AOI22_X1 U2524 ( .A1(VIN), .A2(n3742), .B1(n3720), .B2(n3850), .ZN(
        REGISTER4_n52) );
  AOI22_X1 U2506 ( .A1(VIN), .A2(n3747), .B1(n3705), .B2(n3852), .ZN(
        REGISTER4_n61) );
  AOI22_X1 U2528 ( .A1(VIN), .A2(n3741), .B1(n3675), .B2(n3848), .ZN(
        REGISTER4_n50) );
  AOI22_X1 U2556 ( .A1(VIN), .A2(n3732), .B1(n3695), .B2(n3847), .ZN(
        REGISTER3_n50) );
  AOI22_X1 U2534 ( .A1(VIN), .A2(n3738), .B1(n3704), .B2(n3848), .ZN(
        REGISTER3_n61) );
  AOI22_X1 U2560 ( .A1(VIN), .A2(n3708), .B1(n3761), .B2(n3846), .ZN(
        REGISTER3_n48) );
  AOI22_X1 U2532 ( .A1(VIN), .A2(n3739), .B1(n3773), .B2(n3851), .ZN(
        REGISTER4_n48) );
  AOI22_X1 U2536 ( .A1(VIN), .A2(n3737), .B1(n3700), .B2(n3851), .ZN(
        REGISTER3_n60) );
  AOI22_X1 U2530 ( .A1(VIN), .A2(n3740), .B1(n3706), .B2(n3852), .ZN(
        REGISTER4_n49) );
  NAND2_X1 U2483 ( .A1(VIN), .A2(ff[2]), .ZN(n3250) );
  OAI21_X1 U2482 ( .B1(VIN), .B2(REGISTER_out_n64), .A(n3250), .ZN(
        REGISTER_out_n59) );
  NAND2_X1 U2481 ( .A1(VIN), .A2(ff[1]), .ZN(n3249) );
  OAI21_X1 U2480 ( .B1(VIN), .B2(REGISTER_out_n63), .A(n3249), .ZN(
        REGISTER_out_n60) );
  NAND2_X1 U2479 ( .A1(VIN), .A2(ff[0]), .ZN(n3248) );
  OAI21_X1 U2478 ( .B1(VIN), .B2(REGISTER_out_n62), .A(n3248), .ZN(
        REGISTER_out_n61) );
  NAND2_X1 U2439 ( .A1(n30), .A2(n3848), .ZN(n31) );
  NAND2_X1 U2684 ( .A1(reg2[3]), .A2(VIN), .ZN(n3294) );
  NAND2_X1 U2690 ( .A1(reg2[5]), .A2(VIN), .ZN(n3297) );
  NAND2_X1 U2714 ( .A1(reg2[13]), .A2(VIN), .ZN(n3308) );
  NAND2_X1 U2687 ( .A1(reg2[4]), .A2(VIN), .ZN(n3296) );
  NAND2_X1 U2678 ( .A1(reg2[1]), .A2(VIN), .ZN(n3291) );
  NAND2_X1 U2675 ( .A1(reg2[0]), .A2(VIN), .ZN(n3290) );
  NAND2_X1 U2693 ( .A1(reg2[6]), .A2(VIN), .ZN(n3299) );
  NAND2_X1 U2696 ( .A1(reg2[7]), .A2(VIN), .ZN(n3300) );
  NAND2_X1 U2702 ( .A1(reg2[9]), .A2(VIN), .ZN(n3303) );
  NAND2_X1 U2699 ( .A1(reg2[8]), .A2(VIN), .ZN(n3302) );
  NAND2_X1 U2681 ( .A1(reg2[2]), .A2(VIN), .ZN(n3293) );
  NAND2_X1 U2705 ( .A1(reg2[10]), .A2(VIN), .ZN(n3305) );
  NAND2_X1 U2708 ( .A1(reg2[11]), .A2(VIN), .ZN(n3306) );
  NAND2_X1 U2711 ( .A1(reg2[12]), .A2(VIN), .ZN(n3307) );
  NAND2_X1 U1072 ( .A1(reg2_reg[13]), .A2(n1758), .ZN(n1424) );
  NAND2_X1 U1123 ( .A1(reg2_reg[11]), .A2(n1796), .ZN(n1529) );
  NAND2_X1 U1159 ( .A1(reg2_reg[9]), .A2(n1831), .ZN(n1546) );
  NAND2_X1 U1200 ( .A1(reg2_reg[7]), .A2(n1854), .ZN(n1571) );
  NAND2_X1 U1225 ( .A1(reg2_reg[5]), .A2(n1863), .ZN(n1617) );
  NAND2_X1 U1250 ( .A1(reg2_reg[3]), .A2(n1872), .ZN(n1661) );
  NAND2_X1 U276 ( .A1(reg4_reg[13]), .A2(n859), .ZN(n525) );
  NAND2_X1 U327 ( .A1(reg4_reg[11]), .A2(n897), .ZN(n630) );
  NAND2_X1 U363 ( .A1(reg4_reg[9]), .A2(n932), .ZN(n647) );
  NAND2_X1 U404 ( .A1(reg4_reg[7]), .A2(n955), .ZN(n672) );
  NAND2_X1 U429 ( .A1(reg4_reg[5]), .A2(n964), .ZN(n718) );
  NAND2_X1 U675 ( .A1(reg3_reg[13]), .A2(n1309), .ZN(n975) );
  NAND2_X1 U725 ( .A1(reg3_reg[11]), .A2(n1346), .ZN(n1080) );
  NAND2_X1 U802 ( .A1(reg3_reg[7]), .A2(n1404), .ZN(n1122) );
  NAND2_X1 U761 ( .A1(reg3_reg[9]), .A2(n1381), .ZN(n1097) );
  NAND2_X1 U827 ( .A1(reg3_reg[5]), .A2(n1413), .ZN(n1168) );
  NAND2_X1 U1470 ( .A1(reg1_reg[13]), .A2(n2208), .ZN(n1874) );
  NAND2_X1 U1521 ( .A1(reg1_reg[11]), .A2(n2246), .ZN(n1979) );
  NAND2_X1 U1557 ( .A1(reg1_reg[9]), .A2(n2281), .ZN(n1996) );
  NAND2_X1 U1623 ( .A1(reg1_reg[5]), .A2(n2313), .ZN(n2067) );
  NAND2_X1 U1598 ( .A1(reg1_reg[7]), .A2(n2304), .ZN(n2021) );
  NAND2_X1 U2472 ( .A1(n3235), .A2(n3727), .ZN(n3234) );
  NOR3_X1 U2474 ( .A1(reg7[0]), .A2(reg7[2]), .A3(reg7[1]), .ZN(n3235) );
  NOR2_X1 U2465 ( .A1(reg7[8]), .A2(n3224), .ZN(n3222) );
  NAND2_X1 U679 ( .A1(reg3_reg[11]), .A2(reg3_reg[12]), .ZN(n977) );
  OAI21_X1 U2265 ( .B1(A2[11]), .B2(A2[12]), .A(n2776), .ZN(n3107) );
  NOR2_X1 U2471 ( .A1(reg7[4]), .A2(n3234), .ZN(n3230) );
  NOR2_X1 U2468 ( .A1(reg7[6]), .A2(n3229), .ZN(n3225) );
  NAND2_X1 U1127 ( .A1(reg2_reg[9]), .A2(reg2_reg[10]), .ZN(n1530) );
  NAND2_X1 U331 ( .A1(reg4_reg[9]), .A2(reg4_reg[10]), .ZN(n631) );
  NAND2_X1 U729 ( .A1(reg3_reg[9]), .A2(reg3_reg[10]), .ZN(n1081) );
  NAND2_X1 U2261 ( .A1(A2[13]), .A2(n3107), .ZN(n2774) );
  OAI21_X1 U1874 ( .B1(A1[11]), .B2(A1[12]), .A(n2326), .ZN(n2661) );
  NAND2_X1 U1870 ( .A1(A1[13]), .A2(n2661), .ZN(n2324) );
  NAND2_X1 U1525 ( .A1(reg1_reg[9]), .A2(reg1_reg[10]), .ZN(n1980) );
  NAND2_X1 U1163 ( .A1(reg2_reg[7]), .A2(reg2_reg[8]), .ZN(n1547) );
  NAND2_X1 U367 ( .A1(reg4_reg[7]), .A2(reg4_reg[8]), .ZN(n648) );
  NAND2_X1 U765 ( .A1(reg3_reg[7]), .A2(reg3_reg[8]), .ZN(n1098) );
  NAND2_X1 U1561 ( .A1(reg1_reg[7]), .A2(reg1_reg[8]), .ZN(n1997) );
  OAI21_X1 U2315 ( .B1(A2[9]), .B2(A2[10]), .A(n2880), .ZN(n3144) );
  NAND2_X1 U2311 ( .A1(A2[11]), .A2(n3144), .ZN(n2879) );
  NAND2_X1 U408 ( .A1(reg4_reg[6]), .A2(reg4_reg[5]), .ZN(n673) );
  OAI21_X1 U1924 ( .B1(A1[9]), .B2(A1[10]), .A(n2430), .ZN(n2698) );
  NAND2_X1 U1920 ( .A1(A1[11]), .A2(n2698), .ZN(n2429) );
  INV_X1 U1922 ( .A(A1[11]), .ZN(n2674) );
  OAI21_X1 U1959 ( .B1(A1[7]), .B2(A1[8]), .A(n2447), .ZN(n2733) );
  NAND2_X1 U1955 ( .A1(A1[9]), .A2(n2733), .ZN(n2446) );
  INV_X1 U1957 ( .A(A1[9]), .ZN(n2712) );
  INV_X1 U1696 ( .A(n2445), .ZN(n2435) );
  INV_X1 U1686 ( .A(n2432), .ZN(n2343) );
  INV_X1 U1706 ( .A(n2349), .ZN(n2442) );
  INV_X1 U1700 ( .A(n2350), .ZN(n2443) );
  INV_X1 U2000 ( .A(A1[7]), .ZN(n2409) );
  NAND2_X1 U2021 ( .A1(A1[5]), .A2(n2766), .ZN(n2517) );
  INV_X1 U1732 ( .A(n2494), .ZN(n2477) );
  INV_X1 U1731 ( .A(n2475), .ZN(n2478) );
  INV_X1 U1766 ( .A(n2529), .ZN(n2523) );
  INV_X1 U1744 ( .A(n2511), .ZN(n2486) );
  INV_X1 U1743 ( .A(n2484), .ZN(n2487) );
  INV_X1 U1726 ( .A(n2482), .ZN(n2479) );
  INV_X1 U1725 ( .A(n2483), .ZN(n2480) );
  INV_X1 U1742 ( .A(n2509), .ZN(n2506) );
  INV_X1 U1778 ( .A(n2541), .ZN(n2538) );
  INV_X1 U1777 ( .A(n2542), .ZN(n2540) );
  XOR2_X1 U3178 ( .A(n2549), .B(n2553), .Z(n2550) );
  INV_X1 U1782 ( .A(n2550), .ZN(n2547) );
  INV_X1 U1781 ( .A(n2551), .ZN(n2548) );
  INV_X1 U1784 ( .A(n2546), .ZN(n2543) );
  INV_X1 U1836 ( .A(n2626), .ZN(n2588) );
  INV_X1 U2041 ( .A(A1[0]), .ZN(n2771) );
  INV_X1 U1834 ( .A(n2625), .ZN(n2594) );
  INV_X1 U2031 ( .A(n2337), .ZN(n2335) );
  XOR2_X1 U3195 ( .A(n2619), .B(n2580), .Z(n2581) );
  NOR2_X1 U1802 ( .A1(n2583), .A2(n2381), .ZN(n2378) );
  INV_X1 U1800 ( .A(n2582), .ZN(n2579) );
  INV_X1 U1869 ( .A(n2324), .ZN(n2660) );
  INV_X1 U1919 ( .A(n2429), .ZN(n2697) );
  INV_X1 U1948 ( .A(n2726), .ZN(n2403) );
  INV_X1 U1997 ( .A(n2471), .ZN(n2756) );
  INV_X1 U1979 ( .A(n2334), .ZN(n2339) );
  INV_X1 U1978 ( .A(n2332), .ZN(n2746) );
  INV_X1 U2028 ( .A(n2767), .ZN(n2426) );
  INV_X1 U1972 ( .A(n2405), .ZN(n2739) );
  INV_X1 U1712 ( .A(n2459), .ZN(n2462) );
  INV_X1 U1657 ( .A(n2326), .ZN(n2331) );
  INV_X1 U1076 ( .A(n1431), .ZN(n1426) );
  INV_X1 U1036 ( .A(B1[12]), .ZN(n1425) );
  INV_X1 U1060 ( .A(B1[11]), .ZN(n1534) );
  INV_X1 U1057 ( .A(B1[13]), .ZN(n1430) );
  INV_X1 U888 ( .A(n1532), .ZN(n1443) );
  INV_X1 U1107 ( .A(B1[10]), .ZN(n1541) );
  INV_X1 U898 ( .A(n1545), .ZN(n1535) );
  INV_X1 U908 ( .A(n1449), .ZN(n1542) );
  INV_X1 U1142 ( .A(B1[9]), .ZN(n1553) );
  INV_X1 U1170 ( .A(B1[8]), .ZN(n1555) );
  INV_X1 U902 ( .A(n1450), .ZN(n1543) );
  NAND2_X1 U1204 ( .A1(reg2_reg[6]), .A2(reg2_reg[5]), .ZN(n1572) );
  INV_X1 U1145 ( .A(B1[7]), .ZN(n1567) );
  INV_X1 U914 ( .A(n1559), .ZN(n1562) );
  NAND2_X1 U1229 ( .A1(reg2_reg[3]), .A2(reg2_reg[4]), .ZN(n1618) );
  INV_X1 U928 ( .A(n1582), .ZN(n1579) );
  INV_X1 U927 ( .A(n1583), .ZN(n1580) );
  INV_X1 U934 ( .A(n1594), .ZN(n1577) );
  INV_X1 U1181 ( .A(B1[6]), .ZN(n1591) );
  INV_X1 U933 ( .A(n1575), .ZN(n1578) );
  INV_X1 U968 ( .A(n1629), .ZN(n1623) );
  INV_X1 U1212 ( .A(B1[5]), .ZN(n1613) );
  INV_X1 U946 ( .A(n1611), .ZN(n1586) );
  INV_X1 U945 ( .A(n1584), .ZN(n1587) );
  INV_X1 U944 ( .A(n1609), .ZN(n1606) );
  INV_X1 U980 ( .A(n1641), .ZN(n1638) );
  INV_X1 U979 ( .A(n1642), .ZN(n1640) );
  INV_X1 U1220 ( .A(B1[4]), .ZN(n1625) );
  INV_X1 U984 ( .A(n1650), .ZN(n1647) );
  INV_X1 U983 ( .A(n1651), .ZN(n1648) );
  INV_X1 U1234 ( .A(B1[3]), .ZN(n1665) );
  INV_X1 U986 ( .A(n1646), .ZN(n1643) );
  INV_X1 U1009 ( .A(n1689), .ZN(n1686) );
  INV_X1 U1008 ( .A(n1690), .ZN(n1687) );
  INV_X1 U1027 ( .A(n1703), .ZN(n1702) );
  INV_X1 U1242 ( .A(B1[2]), .ZN(n1683) );
  INV_X1 U1237 ( .A(B1[1]), .ZN(n1436) );
  INV_X1 U1243 ( .A(n1437), .ZN(n1435) );
  INV_X1 U1071 ( .A(n1424), .ZN(n1757) );
  INV_X1 U1231 ( .A(n1864), .ZN(n1526) );
  INV_X1 U1249 ( .A(n1661), .ZN(n1871) );
  INV_X1 U1239 ( .A(n1867), .ZN(n1528) );
  INV_X1 U1224 ( .A(n1617), .ZN(n1862) );
  INV_X1 U1199 ( .A(n1571), .ZN(n1853) );
  INV_X1 U1182 ( .A(n1843), .ZN(n1838) );
  INV_X1 U1194 ( .A(n1512), .ZN(n1851) );
  INV_X1 U1158 ( .A(n1546), .ZN(n1830) );
  INV_X1 U1122 ( .A(n1529), .ZN(n1795) );
  INV_X1 U280 ( .A(n532), .ZN(n527) );
  INV_X1 U240 ( .A(B3[12]), .ZN(n526) );
  INV_X1 U264 ( .A(B3[11]), .ZN(n635) );
  INV_X1 U261 ( .A(B3[13]), .ZN(n531) );
  INV_X1 U92 ( .A(n633), .ZN(n544) );
  INV_X1 U112 ( .A(n550), .ZN(n643) );
  INV_X1 U346 ( .A(B3[9]), .ZN(n654) );
  INV_X1 U374 ( .A(B3[8]), .ZN(n656) );
  INV_X1 U349 ( .A(B3[7]), .ZN(n668) );
  INV_X1 U118 ( .A(n660), .ZN(n663) );
  NAND2_X1 U433 ( .A1(reg4_reg[3]), .A2(reg4_reg[4]), .ZN(n719) );
  INV_X1 U132 ( .A(n683), .ZN(n680) );
  INV_X1 U131 ( .A(n684), .ZN(n681) );
  INV_X1 U138 ( .A(n695), .ZN(n678) );
  INV_X1 U385 ( .A(B3[6]), .ZN(n692) );
  INV_X1 U137 ( .A(n676), .ZN(n679) );
  INV_X1 U184 ( .A(n742), .ZN(n739) );
  INV_X1 U183 ( .A(n743), .ZN(n741) );
  INV_X1 U172 ( .A(n730), .ZN(n724) );
  INV_X1 U424 ( .A(B3[4]), .ZN(n726) );
  INV_X1 U188 ( .A(n751), .ZN(n748) );
  INV_X1 U187 ( .A(n752), .ZN(n749) );
  INV_X1 U438 ( .A(B3[3]), .ZN(n766) );
  INV_X1 U190 ( .A(n747), .ZN(n744) );
  INV_X1 U212 ( .A(n791), .ZN(n788) );
  INV_X1 U231 ( .A(n804), .ZN(n803) );
  INV_X1 U441 ( .A(B3[1]), .ZN(n537) );
  INV_X1 U447 ( .A(n538), .ZN(n536) );
  INV_X1 U435 ( .A(n965), .ZN(n627) );
  INV_X1 U453 ( .A(n762), .ZN(n972) );
  INV_X1 U443 ( .A(n968), .ZN(n629) );
  INV_X1 U428 ( .A(n718), .ZN(n963) );
  INV_X1 U417 ( .A(n950), .ZN(n615) );
  INV_X1 U403 ( .A(n672), .ZN(n954) );
  INV_X1 U386 ( .A(n944), .ZN(n939) );
  INV_X1 U398 ( .A(n613), .ZN(n952) );
  INV_X1 U362 ( .A(n647), .ZN(n931) );
  INV_X1 U356 ( .A(n925), .ZN(n604) );
  INV_X1 U326 ( .A(n630), .ZN(n896) );
  INV_X1 U275 ( .A(n525), .ZN(n858) );
  INV_X1 U150 ( .A(n712), .ZN(n687) );
  INV_X1 U149 ( .A(n685), .ZN(n688) );
  INV_X1 U148 ( .A(n710), .ZN(n707) );
  INV_X1 U102 ( .A(n646), .ZN(n636) );
  INV_X1 U106 ( .A(n551), .ZN(n644) );
  INV_X1 U639 ( .A(B2[12]), .ZN(n976) );
  INV_X1 U660 ( .A(B2[13]), .ZN(n981) );
  INV_X1 U491 ( .A(n1083), .ZN(n994) );
  NAND2_X1 U806 ( .A1(reg3_reg[6]), .A2(reg3_reg[5]), .ZN(n1123) );
  INV_X1 U772 ( .A(B2[8]), .ZN(n1106) );
  INV_X1 U517 ( .A(n1110), .ZN(n1113) );
  INV_X1 U511 ( .A(n1000), .ZN(n1093) );
  INV_X1 U501 ( .A(n1096), .ZN(n1086) );
  NAND2_X1 U831 ( .A1(reg3_reg[3]), .A2(reg3_reg[4]), .ZN(n1169) );
  INV_X1 U531 ( .A(n1133), .ZN(n1130) );
  INV_X1 U530 ( .A(n1134), .ZN(n1131) );
  INV_X1 U537 ( .A(n1145), .ZN(n1128) );
  INV_X1 U536 ( .A(n1126), .ZN(n1129) );
  INV_X1 U571 ( .A(n1180), .ZN(n1174) );
  INV_X1 U549 ( .A(n1162), .ZN(n1137) );
  INV_X1 U548 ( .A(n1135), .ZN(n1138) );
  INV_X1 U547 ( .A(n1160), .ZN(n1157) );
  INV_X1 U583 ( .A(n1192), .ZN(n1189) );
  INV_X1 U582 ( .A(n1193), .ZN(n1191) );
  INV_X1 U822 ( .A(B2[4]), .ZN(n1176) );
  INV_X1 U587 ( .A(n1201), .ZN(n1198) );
  INV_X1 U586 ( .A(n1202), .ZN(n1199) );
  INV_X1 U589 ( .A(n1197), .ZN(n1194) );
  INV_X1 U611 ( .A(n1241), .ZN(n1238) );
  INV_X1 U839 ( .A(B2[1]), .ZN(n987) );
  INV_X1 U845 ( .A(n988), .ZN(n986) );
  INV_X1 U674 ( .A(n975), .ZN(n1308) );
  INV_X1 U833 ( .A(n1414), .ZN(n1077) );
  INV_X1 U851 ( .A(n1212), .ZN(n1421) );
  INV_X1 U841 ( .A(n1417), .ZN(n1079) );
  INV_X1 U826 ( .A(n1168), .ZN(n1412) );
  INV_X1 U815 ( .A(n1399), .ZN(n1065) );
  INV_X1 U801 ( .A(n1122), .ZN(n1403) );
  INV_X1 U784 ( .A(n1393), .ZN(n1388) );
  INV_X1 U796 ( .A(n1063), .ZN(n1401) );
  INV_X1 U760 ( .A(n1097), .ZN(n1380) );
  INV_X1 U724 ( .A(n1080), .ZN(n1345) );
  INV_X1 U505 ( .A(n1001), .ZN(n1094) );
  INV_X1 U1474 ( .A(n1881), .ZN(n1876) );
  INV_X1 U1458 ( .A(B0[11]), .ZN(n1984) );
  INV_X1 U1434 ( .A(B0[12]), .ZN(n1875) );
  INV_X1 U1455 ( .A(B0[13]), .ZN(n1880) );
  INV_X1 U1286 ( .A(n1982), .ZN(n1893) );
  INV_X1 U1296 ( .A(n1995), .ZN(n1985) );
  INV_X1 U1306 ( .A(n1899), .ZN(n1992) );
  INV_X1 U1540 ( .A(B0[9]), .ZN(n2003) );
  NAND2_X1 U1602 ( .A1(reg1_reg[6]), .A2(reg1_reg[5]), .ZN(n2022) );
  NAND2_X1 U1627 ( .A1(reg1_reg[3]), .A2(reg1_reg[4]), .ZN(n2068) );
  INV_X1 U1332 ( .A(n2044), .ZN(n2027) );
  INV_X1 U1331 ( .A(n2025), .ZN(n2028) );
  INV_X1 U1366 ( .A(n2079), .ZN(n2073) );
  INV_X1 U1610 ( .A(B0[5]), .ZN(n2063) );
  INV_X1 U1344 ( .A(n2061), .ZN(n2036) );
  INV_X1 U1343 ( .A(n2034), .ZN(n2037) );
  INV_X1 U1326 ( .A(n2032), .ZN(n2029) );
  INV_X1 U1325 ( .A(n2033), .ZN(n2030) );
  INV_X1 U1342 ( .A(n2059), .ZN(n2056) );
  INV_X1 U1378 ( .A(n2091), .ZN(n2088) );
  INV_X1 U1377 ( .A(n2092), .ZN(n2090) );
  INV_X1 U1618 ( .A(B0[4]), .ZN(n2075) );
  INV_X1 U1382 ( .A(n2100), .ZN(n2097) );
  INV_X1 U1381 ( .A(n2101), .ZN(n2098) );
  INV_X1 U1632 ( .A(B0[3]), .ZN(n2115) );
  INV_X1 U1384 ( .A(n2096), .ZN(n2093) );
  INV_X1 U1406 ( .A(n2140), .ZN(n2137) );
  INV_X1 U1425 ( .A(n2153), .ZN(n2152) );
  INV_X1 U1640 ( .A(B0[2]), .ZN(n2133) );
  INV_X1 U1635 ( .A(B0[1]), .ZN(n1886) );
  INV_X1 U1641 ( .A(n1887), .ZN(n1885) );
  INV_X1 U1469 ( .A(n1874), .ZN(n2207) );
  INV_X1 U1629 ( .A(n2314), .ZN(n1976) );
  INV_X1 U1622 ( .A(n2067), .ZN(n2312) );
  INV_X1 U1611 ( .A(n2299), .ZN(n1964) );
  INV_X1 U1580 ( .A(n2293), .ZN(n2288) );
  INV_X1 U1592 ( .A(n1962), .ZN(n2301) );
  INV_X1 U1550 ( .A(n2274), .ZN(n1953) );
  INV_X1 U1556 ( .A(n1996), .ZN(n2280) );
  INV_X1 U1553 ( .A(n2261), .ZN(n2278) );
  INV_X1 U1520 ( .A(n1979), .ZN(n2245) );
  INV_X1 U1312 ( .A(n2009), .ZN(n2012) );
  INV_X1 U2263 ( .A(A2[13]), .ZN(n2894) );
  INV_X1 U2081 ( .A(n2882), .ZN(n2793) );
  OAI21_X1 U2350 ( .B1(A2[7]), .B2(A2[8]), .A(n2897), .ZN(n3179) );
  NAND2_X1 U2346 ( .A1(A2[9]), .A2(n3179), .ZN(n2896) );
  INV_X1 U2348 ( .A(A2[9]), .ZN(n3158) );
  INV_X1 U2091 ( .A(n2895), .ZN(n2885) );
  INV_X1 U2101 ( .A(n2799), .ZN(n2892) );
  INV_X1 U2095 ( .A(n2800), .ZN(n2893) );
  OAI21_X1 U2393 ( .B1(A2[6]), .B2(A2[5]), .A(n2922), .ZN(n3203) );
  INV_X1 U2391 ( .A(A2[7]), .ZN(n2859) );
  INV_X1 U2438 ( .A(A2[3]), .ZN(n3213) );
  XOR2_X1 U3319 ( .A(n3213), .B(A2[4]), .Z(n3212) );
  NAND2_X1 U2413 ( .A1(A2[5]), .A2(n3212), .ZN(n2967) );
  INV_X1 U2416 ( .A(A2[5]), .ZN(n2873) );
  INV_X1 U2127 ( .A(n2944), .ZN(n2927) );
  INV_X1 U2126 ( .A(n2925), .ZN(n2928) );
  INV_X1 U2161 ( .A(n2982), .ZN(n2973) );
  INV_X1 U2139 ( .A(n2961), .ZN(n2936) );
  INV_X1 U2138 ( .A(n2934), .ZN(n2937) );
  INV_X1 U2121 ( .A(n2932), .ZN(n2929) );
  INV_X1 U2120 ( .A(n2933), .ZN(n2930) );
  INV_X1 U2137 ( .A(n2959), .ZN(n2956) );
  INV_X1 U2171 ( .A(n2990), .ZN(n2987) );
  INV_X1 U2170 ( .A(n2991), .ZN(n2989) );
  INV_X1 U2175 ( .A(n2999), .ZN(n2996) );
  INV_X1 U2174 ( .A(n3000), .ZN(n2997) );
  INV_X1 U2177 ( .A(n2995), .ZN(n2992) );
  INV_X1 U2228 ( .A(n3069), .ZN(n3036) );
  INV_X1 U2431 ( .A(A2[0]), .ZN(n3218) );
  INV_X1 U2226 ( .A(n3068), .ZN(n3042) );
  INV_X1 U2201 ( .A(n3038), .ZN(n3035) );
  INV_X1 U2310 ( .A(n2879), .ZN(n3143) );
  INV_X1 U2421 ( .A(n2787), .ZN(n2785) );
  INV_X1 U2339 ( .A(n3172), .ZN(n2853) );
  INV_X1 U2370 ( .A(n2784), .ZN(n2789) );
  INV_X1 U2369 ( .A(n2782), .ZN(n3192) );
  AND2_X1 U2365 ( .A1(n3188), .A2(n3189), .ZN(n3187) );
  INV_X1 U2418 ( .A(n3214), .ZN(n2876) );
  INV_X1 U2363 ( .A(n2855), .ZN(n3185) );
  INV_X1 U2260 ( .A(n2774), .ZN(n3106) );
  NOR2_X1 U2196 ( .A1(n3031), .A2(n2831), .ZN(n2827) );
  INV_X1 U2195 ( .A(n3030), .ZN(n3027) );
  INV_X1 U2107 ( .A(n2909), .ZN(n2912) );
  INV_X1 U2049 ( .A(p10_final_product2_26_), .ZN(p10_final_product2_25_) );
  INV_X1 U2052 ( .A(n2776), .ZN(n2781) );
  INV_X1 U2441 ( .A(n3222), .ZN(n3221) );
  INV_X1 U2445 ( .A(n3225), .ZN(n3228) );
  INV_X1 U2449 ( .A(n3230), .ZN(n3233) );
  INV_X1 U2453 ( .A(n3235), .ZN(n3238) );
  INV_X1 U2522 ( .A(n3270), .ZN(REGISTER4_n53) );
  INV_X1 U2514 ( .A(n3266), .ZN(REGISTER4_n57) );
  INV_X1 U2546 ( .A(n3282), .ZN(REGISTER3_n55) );
  INV_X1 U2518 ( .A(n3268), .ZN(REGISTER4_n55) );
  INV_X1 U2558 ( .A(n3288), .ZN(REGISTER3_n49) );
  INV_X1 U2538 ( .A(n3278), .ZN(REGISTER3_n59) );
  INV_X1 U2554 ( .A(n3286), .ZN(REGISTER3_n51) );
  INV_X1 U2542 ( .A(n3280), .ZN(REGISTER3_n57) );
  INV_X1 U2510 ( .A(n3264), .ZN(REGISTER4_n59) );
  INV_X1 U2550 ( .A(n3284), .ZN(REGISTER3_n53) );
  DFFR_X2 REGISTER1_q_reg_1_ ( .D(REGISTER1_n60), .CK(CLK), .RN(RST_n), .Q(
        reg1_reg[1]), .QN(n3715) );
  OR2_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U1 ( .A1(n3466), .A2(reg7[0]), 
        .ZN(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_) );
  XNOR2_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2 ( .A(reg7[0]), .B(n3466), 
        .ZN(fb_0_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_1 ( .A(SUB1_N1), .B(n3474), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_1_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_), .S(fb_1_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_2 ( .A(SUB1_N2), .B(n3473), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_2_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_), .S(fb_2_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_3 ( .A(SUB1_N3), .B(n3472), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_3_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_), .S(fb_3_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_4 ( .A(SUB1_N4), .B(n3471), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_4_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_), .S(fb_4_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_5 ( .A(SUB1_N5), .B(n3470), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_5_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_), .S(fb_5_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_6 ( .A(SUB1_N6), .B(n3469), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_6_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_), .S(fb_6_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_7 ( .A(SUB1_N7), .B(n3468), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_7_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_), .S(fb_7_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_8 ( .A(SUB1_N8), .B(n3467), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_8_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_), .S(fb_8_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_9 ( .A(SUB1_N9), .B(n3479), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_9_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_), .S(fb_9_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_10 ( .A(SUB1_N10), .B(n3478), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_10_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_), .S(fb_10_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_11 ( .A(SUB1_N11), .B(n3477), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_11_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_), .S(fb_11_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_12 ( .A(SUB1_N12), .B(n3476), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_12_), .CO(
        SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_), .S(fb_12_) );
  FA_X1 SUB1_sub_0_root_sub_0_root_sub_21_2_U2_13 ( .A(SUB1_N13), .B(n3475), 
        .CI(SUB1_sub_0_root_sub_0_root_sub_21_2_carry_13_), .S(fb_13_) );
  AND2_X1 s6_add_23_U1 ( .A1(mul1_reg[0]), .A2(mul2_reg[0]), .ZN(
        s6_add_23_carry_1_) );
  XOR2_X1 s6_add_23_U2 ( .A(mul2_reg[0]), .B(mul1_reg[0]), .Z(sig_ff1_0_) );
  FA_X1 s6_add_23_U1_1 ( .A(mul1_reg[1]), .B(mul2_reg[1]), .CI(
        s6_add_23_carry_1_), .CO(s6_add_23_carry_2_), .S(sig_ff1_1_) );
  FA_X1 s6_add_23_U1_2 ( .A(mul1_reg[2]), .B(mul2_reg[2]), .CI(
        s6_add_23_carry_2_), .CO(s6_add_23_carry_3_), .S(sig_ff1_2_) );
  FA_X1 s6_add_23_U1_3 ( .A(mul1_reg[3]), .B(mul2_reg[3]), .CI(
        s6_add_23_carry_3_), .CO(s6_add_23_carry_4_), .S(sig_ff1_3_) );
  FA_X1 s6_add_23_U1_4 ( .A(mul1_reg[4]), .B(mul2_reg[4]), .CI(
        s6_add_23_carry_4_), .CO(s6_add_23_carry_5_), .S(sig_ff1_4_) );
  FA_X1 s6_add_23_U1_5 ( .A(mul1_reg[5]), .B(mul2_reg[5]), .CI(
        s6_add_23_carry_5_), .CO(s6_add_23_carry_6_), .S(sig_ff1_5_) );
  FA_X1 s6_add_23_U1_6 ( .A(mul1_reg[6]), .B(mul2_reg[6]), .CI(
        s6_add_23_carry_6_), .CO(s6_add_23_carry_7_), .S(sig_ff1_6_) );
  FA_X1 s6_add_23_U1_7 ( .A(mul1_reg[7]), .B(mul2_reg[7]), .CI(
        s6_add_23_carry_7_), .CO(s6_add_23_carry_8_), .S(sig_ff1_7_) );
  FA_X1 s6_add_23_U1_8 ( .A(mul1_reg[8]), .B(mul2_reg[8]), .CI(
        s6_add_23_carry_8_), .CO(s6_add_23_carry_9_), .S(sig_ff1_8_) );
  FA_X1 s6_add_23_U1_9 ( .A(mul1_reg[9]), .B(mul2_reg[9]), .CI(
        s6_add_23_carry_9_), .CO(s6_add_23_carry_10_), .S(sig_ff1_9_) );
  FA_X1 s6_add_23_U1_10 ( .A(mul1_reg[10]), .B(mul2_reg[10]), .CI(
        s6_add_23_carry_10_), .CO(s6_add_23_carry_11_), .S(sig_ff1_10_) );
  FA_X1 s6_add_23_U1_11 ( .A(mul1_reg[11]), .B(mul2_reg[11]), .CI(
        s6_add_23_carry_11_), .CO(s6_add_23_carry_12_), .S(sig_ff1_11_) );
  FA_X1 s6_add_23_U1_12 ( .A(mul1_reg[12]), .B(mul2_reg[12]), .CI(
        s6_add_23_carry_12_), .CO(s6_add_23_carry_13_), .S(sig_ff1_12_) );
  FA_X1 s6_add_23_U1_13 ( .A(mul1_reg[13]), .B(mul2_reg[13]), .CI(
        s6_add_23_carry_13_), .S(sig_ff1_13_) );
  AND2_X1 s9_add_23_U1 ( .A1(fb_0_), .A2(xin[0]), .ZN(s9_add_23_carry_1_) );
  FA_X1 s9_add_23_U1_1 ( .A(fb_1_), .B(xin[1]), .CI(s9_add_23_carry_1_), .CO(
        s9_add_23_carry_2_), .S(w[1]) );
  FA_X1 s9_add_23_U1_2 ( .A(fb_2_), .B(xin[2]), .CI(s9_add_23_carry_2_), .CO(
        s9_add_23_carry_3_), .S(w[2]) );
  FA_X1 s9_add_23_U1_3 ( .A(fb_3_), .B(xin[3]), .CI(s9_add_23_carry_3_), .CO(
        s9_add_23_carry_4_), .S(w[3]) );
  FA_X1 s9_add_23_U1_4 ( .A(fb_4_), .B(xin[4]), .CI(s9_add_23_carry_4_), .CO(
        s9_add_23_carry_5_), .S(w[4]) );
  FA_X1 s9_add_23_U1_5 ( .A(fb_5_), .B(xin[5]), .CI(s9_add_23_carry_5_), .CO(
        s9_add_23_carry_6_), .S(w[5]) );
  FA_X1 s9_add_23_U1_6 ( .A(fb_6_), .B(xin[6]), .CI(s9_add_23_carry_6_), .CO(
        s9_add_23_carry_7_), .S(w[6]) );
  FA_X1 s9_add_23_U1_7 ( .A(fb_7_), .B(xin[7]), .CI(s9_add_23_carry_7_), .CO(
        s9_add_23_carry_8_), .S(w[7]) );
  FA_X1 s9_add_23_U1_8 ( .A(fb_8_), .B(xin[8]), .CI(s9_add_23_carry_8_), .CO(
        s9_add_23_carry_9_), .S(w[8]) );
  FA_X1 s9_add_23_U1_9 ( .A(fb_9_), .B(xin[9]), .CI(s9_add_23_carry_9_), .CO(
        s9_add_23_carry_10_), .S(w[9]) );
  FA_X1 s9_add_23_U1_10 ( .A(fb_10_), .B(xin[10]), .CI(s9_add_23_carry_10_), 
        .CO(s9_add_23_carry_11_), .S(w[10]) );
  FA_X1 s9_add_23_U1_11 ( .A(fb_11_), .B(xin[11]), .CI(s9_add_23_carry_11_), 
        .CO(s9_add_23_carry_12_), .S(w[11]) );
  FA_X1 s9_add_23_U1_12 ( .A(fb_12_), .B(xin[12]), .CI(s9_add_23_carry_12_), 
        .CO(s9_add_23_carry_13_), .S(w[12]) );
  FA_X1 s9_add_23_U1_13 ( .A(fb_13_), .B(xin[13]), .CI(s9_add_23_carry_13_), 
        .S(w[13]) );
  AND2_X1 s8_add_23_U1 ( .A1(sig_ff1_0_), .A2(sig_ff2_0_), .ZN(
        s8_add_23_carry_1_) );
  XOR2_X1 s8_add_23_U2 ( .A(sig_ff2_0_), .B(sig_ff1_0_), .Z(ff[0]) );
  FA_X1 s8_add_23_U1_1 ( .A(sig_ff1_1_), .B(sig_ff2_1_), .CI(
        s8_add_23_carry_1_), .CO(s8_add_23_carry_2_), .S(ff[1]) );
  FA_X1 s8_add_23_U1_2 ( .A(sig_ff1_2_), .B(sig_ff2_2_), .CI(
        s8_add_23_carry_2_), .CO(s8_add_23_carry_3_), .S(ff[2]) );
  FA_X1 s8_add_23_U1_3 ( .A(sig_ff1_3_), .B(sig_ff2_3_), .CI(
        s8_add_23_carry_3_), .CO(s8_add_23_carry_4_), .S(ff[3]) );
  FA_X1 s8_add_23_U1_4 ( .A(sig_ff1_4_), .B(sig_ff2_4_), .CI(
        s8_add_23_carry_4_), .CO(s8_add_23_carry_5_), .S(ff[4]) );
  FA_X1 s8_add_23_U1_5 ( .A(sig_ff1_5_), .B(sig_ff2_5_), .CI(
        s8_add_23_carry_5_), .CO(s8_add_23_carry_6_), .S(ff[5]) );
  FA_X1 s8_add_23_U1_6 ( .A(sig_ff1_6_), .B(sig_ff2_6_), .CI(
        s8_add_23_carry_6_), .CO(s8_add_23_carry_7_), .S(ff[6]) );
  FA_X1 s8_add_23_U1_7 ( .A(sig_ff1_7_), .B(sig_ff2_7_), .CI(
        s8_add_23_carry_7_), .CO(s8_add_23_carry_8_), .S(ff[7]) );
  FA_X1 s8_add_23_U1_8 ( .A(sig_ff1_8_), .B(sig_ff2_8_), .CI(
        s8_add_23_carry_8_), .CO(s8_add_23_carry_9_), .S(ff[8]) );
  FA_X1 s8_add_23_U1_9 ( .A(sig_ff1_9_), .B(sig_ff2_9_), .CI(
        s8_add_23_carry_9_), .CO(s8_add_23_carry_10_), .S(ff[9]) );
  FA_X1 s8_add_23_U1_10 ( .A(sig_ff1_10_), .B(sig_ff2_10_), .CI(
        s8_add_23_carry_10_), .CO(s8_add_23_carry_11_), .S(ff[10]) );
  FA_X1 s8_add_23_U1_11 ( .A(sig_ff1_11_), .B(sig_ff2_11_), .CI(
        s8_add_23_carry_11_), .CO(s8_add_23_carry_12_), .S(ff[11]) );
  FA_X1 s8_add_23_U1_12 ( .A(sig_ff1_12_), .B(sig_ff2_12_), .CI(
        s8_add_23_carry_12_), .CO(s8_add_23_carry_13_), .S(ff[12]) );
  FA_X1 s8_add_23_U1_13 ( .A(sig_ff1_13_), .B(sig_ff2_13_), .CI(
        s8_add_23_carry_13_), .S(ff[13]) );
  AND2_X1 s7_add_23_U1 ( .A1(mul3_reg[0]), .A2(mul4_reg[0]), .ZN(
        s7_add_23_carry_1_) );
  XOR2_X1 s7_add_23_U2 ( .A(mul4_reg[0]), .B(mul3_reg[0]), .Z(sig_ff2_0_) );
  FA_X1 s7_add_23_U1_1 ( .A(mul3_reg[1]), .B(mul4_reg[1]), .CI(
        s7_add_23_carry_1_), .CO(s7_add_23_carry_2_), .S(sig_ff2_1_) );
  FA_X1 s7_add_23_U1_2 ( .A(mul3_reg[2]), .B(mul4_reg[2]), .CI(
        s7_add_23_carry_2_), .CO(s7_add_23_carry_3_), .S(sig_ff2_2_) );
  FA_X1 s7_add_23_U1_3 ( .A(mul3_reg[3]), .B(mul4_reg[3]), .CI(
        s7_add_23_carry_3_), .CO(s7_add_23_carry_4_), .S(sig_ff2_3_) );
  FA_X1 s7_add_23_U1_4 ( .A(mul3_reg[4]), .B(mul4_reg[4]), .CI(
        s7_add_23_carry_4_), .CO(s7_add_23_carry_5_), .S(sig_ff2_4_) );
  FA_X1 s7_add_23_U1_5 ( .A(mul3_reg[5]), .B(mul4_reg[5]), .CI(
        s7_add_23_carry_5_), .CO(s7_add_23_carry_6_), .S(sig_ff2_5_) );
  FA_X1 s7_add_23_U1_6 ( .A(mul3_reg[6]), .B(mul4_reg[6]), .CI(
        s7_add_23_carry_6_), .CO(s7_add_23_carry_7_), .S(sig_ff2_6_) );
  FA_X1 s7_add_23_U1_7 ( .A(mul3_reg[7]), .B(mul4_reg[7]), .CI(
        s7_add_23_carry_7_), .CO(s7_add_23_carry_8_), .S(sig_ff2_7_) );
  FA_X1 s7_add_23_U1_8 ( .A(mul3_reg[8]), .B(mul4_reg[8]), .CI(
        s7_add_23_carry_8_), .CO(s7_add_23_carry_9_), .S(sig_ff2_8_) );
  FA_X1 s7_add_23_U1_9 ( .A(mul3_reg[9]), .B(mul4_reg[9]), .CI(
        s7_add_23_carry_9_), .CO(s7_add_23_carry_10_), .S(sig_ff2_9_) );
  FA_X1 s7_add_23_U1_10 ( .A(mul3_reg[10]), .B(mul4_reg[10]), .CI(
        s7_add_23_carry_10_), .CO(s7_add_23_carry_11_), .S(sig_ff2_10_) );
  FA_X1 s7_add_23_U1_11 ( .A(mul3_reg[11]), .B(mul4_reg[11]), .CI(
        s7_add_23_carry_11_), .CO(s7_add_23_carry_12_), .S(sig_ff2_11_) );
  FA_X1 s7_add_23_U1_12 ( .A(mul3_reg[12]), .B(mul4_reg[12]), .CI(
        s7_add_23_carry_12_), .CO(s7_add_23_carry_13_), .S(sig_ff2_12_) );
  FA_X1 s7_add_23_U1_13 ( .A(mul3_reg[13]), .B(mul4_reg[13]), .CI(
        s7_add_23_carry_13_), .S(sig_ff2_13_) );
  INV_X1 p6_Partial_products_sum_add_23_U40 ( .A(p6_C[53]), .ZN(
        p6_Partial_products_sum_add_23_n178) );
  INV_X1 p6_Partial_products_sum_add_23_U39 ( .A(p6_S[54]), .ZN(
        p6_Partial_products_sum_add_23_n177) );
  INV_X1 p6_Partial_products_sum_add_23_U48 ( .A(p6_C[51]), .ZN(
        p6_Partial_products_sum_add_23_n184) );
  INV_X1 p6_Partial_products_sum_add_23_U47 ( .A(p6_S[52]), .ZN(
        p6_Partial_products_sum_add_23_n183) );
  INV_X1 p6_Partial_products_sum_add_23_U64 ( .A(p6_C[47]), .ZN(
        p6_Partial_products_sum_add_23_n196) );
  INV_X1 p6_Partial_products_sum_add_23_U63 ( .A(p6_S[48]), .ZN(
        p6_Partial_products_sum_add_23_n195) );
  INV_X1 p6_Partial_products_sum_add_23_U72 ( .A(p6_C[45]), .ZN(
        p6_Partial_products_sum_add_23_n202) );
  INV_X1 p6_Partial_products_sum_add_23_U71 ( .A(p6_S[46]), .ZN(
        p6_Partial_products_sum_add_23_n201) );
  INV_X1 p6_Partial_products_sum_add_23_U80 ( .A(p6_C[43]), .ZN(
        p6_Partial_products_sum_add_23_n208) );
  INV_X1 p6_Partial_products_sum_add_23_U79 ( .A(p6_S[44]), .ZN(
        p6_Partial_products_sum_add_23_n207) );
  INV_X1 p6_Partial_products_sum_add_23_U55 ( .A(p6_S[50]), .ZN(
        p6_Partial_products_sum_add_23_n189) );
  INV_X1 p6_Partial_products_sum_add_23_U56 ( .A(p6_C[49]), .ZN(
        p6_Partial_products_sum_add_23_n190) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U82 ( .A(
        p6_Partial_products_sum_add_23_n211), .B(
        p6_Partial_products_sum_add_23_n210), .ZN(temp1[0]) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U109 ( .A(p6_S[43]), .B(p6_C[42]), 
        .ZN(p6_Partial_products_sum_add_23_n211) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U77 ( .A(
        p6_Partial_products_sum_add_23_n206), .B(
        p6_Partial_products_sum_add_23_n209), .ZN(temp1[1]) );
  AOI22_X1 p6_Partial_products_sum_add_23_U78 ( .A1(p6_S[44]), .A2(p6_C[43]), 
        .B1(p6_Partial_products_sum_add_23_n208), .B2(
        p6_Partial_products_sum_add_23_n207), .ZN(
        p6_Partial_products_sum_add_23_n209) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U74 ( .A(
        p6_Partial_products_sum_add_23_n205), .B(
        p6_Partial_products_sum_add_23_n204), .ZN(temp1[2]) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U76 ( .A(p6_S[45]), .B(p6_C[44]), 
        .ZN(p6_Partial_products_sum_add_23_n205) );
  AOI22_X1 p6_Partial_products_sum_add_23_U70 ( .A1(p6_S[46]), .A2(p6_C[45]), 
        .B1(p6_Partial_products_sum_add_23_n202), .B2(
        p6_Partial_products_sum_add_23_n201), .ZN(
        p6_Partial_products_sum_add_23_n203) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U68 ( .A(p6_S[47]), .B(p6_C[46]), 
        .ZN(p6_Partial_products_sum_add_23_n199) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U61 ( .A(
        p6_Partial_products_sum_add_23_n194), .B(
        p6_Partial_products_sum_add_23_n197), .ZN(temp1[5]) );
  AOI22_X1 p6_Partial_products_sum_add_23_U62 ( .A1(p6_S[48]), .A2(p6_C[47]), 
        .B1(p6_Partial_products_sum_add_23_n196), .B2(
        p6_Partial_products_sum_add_23_n195), .ZN(
        p6_Partial_products_sum_add_23_n197) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U60 ( .A(p6_S[49]), .B(p6_C[48]), 
        .ZN(p6_Partial_products_sum_add_23_n193) );
  AOI22_X1 p6_Partial_products_sum_add_23_U54 ( .A1(p6_S[50]), .A2(p6_C[49]), 
        .B1(p6_Partial_products_sum_add_23_n190), .B2(
        p6_Partial_products_sum_add_23_n189), .ZN(
        p6_Partial_products_sum_add_23_n191) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U52 ( .A(p6_S[51]), .B(p6_C[50]), 
        .ZN(p6_Partial_products_sum_add_23_n187) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U45 ( .A(
        p6_Partial_products_sum_add_23_n182), .B(
        p6_Partial_products_sum_add_23_n185), .ZN(temp1[9]) );
  AOI22_X1 p6_Partial_products_sum_add_23_U46 ( .A1(p6_S[52]), .A2(p6_C[51]), 
        .B1(p6_Partial_products_sum_add_23_n184), .B2(
        p6_Partial_products_sum_add_23_n183), .ZN(
        p6_Partial_products_sum_add_23_n185) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U44 ( .A(p6_S[53]), .B(p6_C[52]), 
        .ZN(p6_Partial_products_sum_add_23_n181) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U37 ( .A(
        p6_Partial_products_sum_add_23_n176), .B(
        p6_Partial_products_sum_add_23_n179), .ZN(temp1[11]) );
  AOI22_X1 p6_Partial_products_sum_add_23_U38 ( .A1(p6_S[54]), .A2(p6_C[53]), 
        .B1(p6_Partial_products_sum_add_23_n178), .B2(
        p6_Partial_products_sum_add_23_n177), .ZN(
        p6_Partial_products_sum_add_23_n179) );
  XNOR2_X1 p6_Partial_products_sum_add_23_U36 ( .A(p6_C[54]), .B(
        p6_final_product2_25_), .ZN(p6_Partial_products_sum_add_23_n175) );
  NAND2_X1 p6_Partial_products_sum_add_23_U88 ( .A1(p6_C[39]), .A2(p6_S[40]), 
        .ZN(p6_Partial_products_sum_add_23_n218) );
  NOR2_X1 p6_Partial_products_sum_add_23_U89 ( .A1(p6_C[39]), .A2(p6_S[40]), 
        .ZN(p6_Partial_products_sum_add_23_n217) );
  NAND2_X1 p6_Partial_products_sum_add_23_U92 ( .A1(p6_C[37]), .A2(p6_S[38]), 
        .ZN(p6_Partial_products_sum_add_23_n222) );
  NOR2_X1 p6_Partial_products_sum_add_23_U93 ( .A1(p6_C[37]), .A2(p6_S[38]), 
        .ZN(p6_Partial_products_sum_add_23_n221) );
  NAND2_X1 p6_Partial_products_sum_add_23_U96 ( .A1(p6_C[35]), .A2(p6_S[36]), 
        .ZN(p6_Partial_products_sum_add_23_n226) );
  NOR2_X1 p6_Partial_products_sum_add_23_U97 ( .A1(p6_C[35]), .A2(p6_S[36]), 
        .ZN(p6_Partial_products_sum_add_23_n225) );
  NAND2_X1 p6_Partial_products_sum_add_23_U100 ( .A1(p6_S[34]), .A2(p6_C[33]), 
        .ZN(p6_Partial_products_sum_add_23_n230) );
  NOR2_X1 p6_Partial_products_sum_add_23_U101 ( .A1(p6_S[34]), .A2(p6_C[33]), 
        .ZN(p6_Partial_products_sum_add_23_n229) );
  NAND2_X1 p6_Partial_products_sum_add_23_U104 ( .A1(n3654), .A2(reg1_reg[3]), 
        .ZN(p6_Partial_products_sum_add_23_n233) );
  INV_X1 p10_Partial_products_sum_add_23_U53 ( .A(p10_C[51]), .ZN(
        p10_Partial_products_sum_add_23_n291) );
  INV_X1 p10_Partial_products_sum_add_23_U52 ( .A(p10_S[52]), .ZN(
        p10_Partial_products_sum_add_23_n290) );
  INV_X1 p10_Partial_products_sum_add_23_U77 ( .A(p10_C[45]), .ZN(
        p10_Partial_products_sum_add_23_n309) );
  INV_X1 p10_Partial_products_sum_add_23_U76 ( .A(p10_S[46]), .ZN(
        p10_Partial_products_sum_add_23_n308) );
  INV_X1 p10_Partial_products_sum_add_23_U85 ( .A(p10_C[43]), .ZN(
        p10_Partial_products_sum_add_23_n315) );
  INV_X1 p10_Partial_products_sum_add_23_U84 ( .A(p10_S[44]), .ZN(
        p10_Partial_products_sum_add_23_n314) );
  INV_X1 p10_Partial_products_sum_add_23_U69 ( .A(p10_C[47]), .ZN(
        p10_Partial_products_sum_add_23_n303) );
  INV_X1 p10_Partial_products_sum_add_23_U60 ( .A(p10_S[50]), .ZN(
        p10_Partial_products_sum_add_23_n296) );
  INV_X1 p10_Partial_products_sum_add_23_U61 ( .A(p10_C[49]), .ZN(
        p10_Partial_products_sum_add_23_n297) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U115 ( .A(p10_S[43]), .B(p10_C[42]), 
        .ZN(p10_Partial_products_sum_add_23_n318) );
  AOI22_X1 p10_Partial_products_sum_add_23_U83 ( .A1(p10_S[44]), .A2(p10_C[43]), .B1(p10_Partial_products_sum_add_23_n315), .B2(
        p10_Partial_products_sum_add_23_n314), .ZN(
        p10_Partial_products_sum_add_23_n316) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U81 ( .A(p10_S[45]), .B(p10_C[44]), 
        .ZN(p10_Partial_products_sum_add_23_n312) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U74 ( .A(
        p10_Partial_products_sum_add_23_n307), .B(
        p10_Partial_products_sum_add_23_n310), .ZN(temp5[3]) );
  AOI22_X1 p10_Partial_products_sum_add_23_U75 ( .A1(p10_S[46]), .A2(p10_C[45]), .B1(p10_Partial_products_sum_add_23_n309), .B2(
        p10_Partial_products_sum_add_23_n308), .ZN(
        p10_Partial_products_sum_add_23_n310) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U73 ( .A(p10_S[47]), .B(p10_C[46]), 
        .ZN(p10_Partial_products_sum_add_23_n306) );
  AOI22_X1 p10_Partial_products_sum_add_23_U67 ( .A1(p10_S[48]), .A2(p10_C[47]), .B1(p10_Partial_products_sum_add_23_n303), .B2(
        p10_Partial_products_sum_add_23_n302), .ZN(
        p10_Partial_products_sum_add_23_n304) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U65 ( .A(p10_S[49]), .B(p10_C[48]), 
        .ZN(p10_Partial_products_sum_add_23_n300) );
  AOI22_X1 p10_Partial_products_sum_add_23_U59 ( .A1(p10_S[50]), .A2(p10_C[49]), .B1(p10_Partial_products_sum_add_23_n297), .B2(
        p10_Partial_products_sum_add_23_n296), .ZN(
        p10_Partial_products_sum_add_23_n298) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U57 ( .A(p10_S[51]), .B(p10_C[50]), 
        .ZN(p10_Partial_products_sum_add_23_n294) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U50 ( .A(
        p10_Partial_products_sum_add_23_n289), .B(
        p10_Partial_products_sum_add_23_n292), .ZN(temp5[9]) );
  AOI22_X1 p10_Partial_products_sum_add_23_U51 ( .A1(p10_S[52]), .A2(p10_C[51]), .B1(p10_Partial_products_sum_add_23_n291), .B2(
        p10_Partial_products_sum_add_23_n290), .ZN(
        p10_Partial_products_sum_add_23_n292) );
  XNOR2_X1 p10_Partial_products_sum_add_23_U49 ( .A(p10_S[53]), .B(p10_C[52]), 
        .ZN(p10_Partial_products_sum_add_23_n288) );
  AOI22_X1 p10_Partial_products_sum_add_23_U42 ( .A1(p10_C[53]), .A2(p10_S[54]), .B1(p10_Partial_products_sum_add_23_n285), .B2(
        p10_Partial_products_sum_add_23_n284), .ZN(
        p10_Partial_products_sum_add_23_n286) );
  AOI22_X1 p10_Partial_products_sum_add_23_U38 ( .A1(p10_final_product2_25_), 
        .A2(p10_Partial_products_sum_add_23_n277), .B1(p10_C[54]), .B2(
        p10_final_product2_26_), .ZN(p10_Partial_products_sum_add_23_n281) );
  NAND2_X1 p10_Partial_products_sum_add_23_U97 ( .A1(
        p10_Partial_products_sum_add_23_n329), .A2(p10_S[38]), .ZN(
        p10_Partial_products_sum_add_23_n328) );
  OAI21_X1 p10_Partial_products_sum_add_23_U98 ( .B1(
        p10_Partial_products_sum_add_23_n329), .B2(p10_S[38]), .A(p10_C[37]), 
        .ZN(p10_Partial_products_sum_add_23_n327) );
  NAND2_X1 p10_Partial_products_sum_add_23_U99 ( .A1(
        p10_Partial_products_sum_add_23_n330), .A2(
        p10_Partial_products_sum_add_23_n331), .ZN(
        p10_Partial_products_sum_add_23_n329) );
  NAND2_X1 p10_Partial_products_sum_add_23_U100 ( .A1(p10_S[37]), .A2(
        p10_C[36]), .ZN(p10_Partial_products_sum_add_23_n331) );
  OAI21_X1 p10_Partial_products_sum_add_23_U101 ( .B1(p10_S[37]), .B2(
        p10_C[36]), .A(p10_Partial_products_sum_add_23_n332), .ZN(
        p10_Partial_products_sum_add_23_n330) );
  NAND2_X1 p10_Partial_products_sum_add_23_U103 ( .A1(p10_C[35]), .A2(
        p10_S[36]), .ZN(p10_Partial_products_sum_add_23_n335) );
  NOR2_X1 p10_Partial_products_sum_add_23_U104 ( .A1(p10_C[35]), .A2(p10_S[36]), .ZN(p10_Partial_products_sum_add_23_n334) );
  NAND2_X1 p10_Partial_products_sum_add_23_U107 ( .A1(p10_C[33]), .A2(
        p10_S[34]), .ZN(p10_Partial_products_sum_add_23_n339) );
  XOR2_X1 p10_Partial_products_sum_add_23_U116 ( .A(
        p10_Partial_products_sum_add_23_n280), .B(
        p10_Partial_products_sum_add_23_n286), .Z(temp5[11]) );
  INV_X1 p11_Partial_products_sum_add_23_U48 ( .A(p11_C[51]), .ZN(
        p11_Partial_products_sum_add_23_n267) );
  INV_X1 p11_Partial_products_sum_add_23_U47 ( .A(p11_S[52]), .ZN(
        p11_Partial_products_sum_add_23_n266) );
  INV_X1 p11_Partial_products_sum_add_23_U64 ( .A(p11_C[47]), .ZN(
        p11_Partial_products_sum_add_23_n279) );
  INV_X1 p11_Partial_products_sum_add_23_U63 ( .A(p11_S[48]), .ZN(
        p11_Partial_products_sum_add_23_n278) );
  INV_X1 p11_Partial_products_sum_add_23_U72 ( .A(p11_C[45]), .ZN(
        p11_Partial_products_sum_add_23_n285) );
  INV_X1 p11_Partial_products_sum_add_23_U71 ( .A(p11_S[46]), .ZN(
        p11_Partial_products_sum_add_23_n284) );
  AND2_X1 p11_Partial_products_sum_add_23_U107 ( .A1(A1[1]), .A2(
        p11_final_product1[0]), .ZN(p11_Partial_products_sum_add_23_n318) );
  INV_X1 p11_Partial_products_sum_add_23_U55 ( .A(p11_S[50]), .ZN(
        p11_Partial_products_sum_add_23_n272) );
  INV_X1 p11_Partial_products_sum_add_23_U56 ( .A(p11_C[49]), .ZN(
        p11_Partial_products_sum_add_23_n273) );
  INV_X1 p11_Partial_products_sum_add_23_U39 ( .A(p11_S[54]), .ZN(
        p11_Partial_products_sum_add_23_n260) );
  INV_X1 p11_Partial_products_sum_add_23_U40 ( .A(p11_C[53]), .ZN(
        p11_Partial_products_sum_add_23_n261) );
  XNOR2_X1 p11_Partial_products_sum_add_23_U76 ( .A(p11_S[45]), .B(p11_C[44]), 
        .ZN(p11_Partial_products_sum_add_23_n288) );
  AOI22_X1 p11_Partial_products_sum_add_23_U70 ( .A1(p11_S[46]), .A2(p11_C[45]), .B1(p11_Partial_products_sum_add_23_n285), .B2(
        p11_Partial_products_sum_add_23_n284), .ZN(
        p11_Partial_products_sum_add_23_n286) );
  AOI22_X1 p11_Partial_products_sum_add_23_U62 ( .A1(p11_S[48]), .A2(p11_C[47]), .B1(p11_Partial_products_sum_add_23_n279), .B2(
        p11_Partial_products_sum_add_23_n278), .ZN(
        p11_Partial_products_sum_add_23_n280) );
  XNOR2_X1 p11_Partial_products_sum_add_23_U60 ( .A(p11_S[49]), .B(p11_C[48]), 
        .ZN(p11_Partial_products_sum_add_23_n276) );
  AOI22_X1 p11_Partial_products_sum_add_23_U54 ( .A1(p11_S[50]), .A2(p11_C[49]), .B1(p11_Partial_products_sum_add_23_n273), .B2(
        p11_Partial_products_sum_add_23_n272), .ZN(
        p11_Partial_products_sum_add_23_n274) );
  XNOR2_X1 p11_Partial_products_sum_add_23_U52 ( .A(p11_S[51]), .B(p11_C[50]), 
        .ZN(p11_Partial_products_sum_add_23_n270) );
  AOI22_X1 p11_Partial_products_sum_add_23_U46 ( .A1(p11_S[52]), .A2(p11_C[51]), .B1(p11_Partial_products_sum_add_23_n267), .B2(
        p11_Partial_products_sum_add_23_n266), .ZN(
        p11_Partial_products_sum_add_23_n268) );
  XNOR2_X1 p11_Partial_products_sum_add_23_U44 ( .A(p11_S[53]), .B(p11_C[52]), 
        .ZN(p11_Partial_products_sum_add_23_n264) );
  AOI22_X1 p11_Partial_products_sum_add_23_U38 ( .A1(p11_S[54]), .A2(p11_C[53]), .B1(p11_Partial_products_sum_add_23_n261), .B2(
        p11_Partial_products_sum_add_23_n260), .ZN(
        p11_Partial_products_sum_add_23_n262) );
  XNOR2_X1 p11_Partial_products_sum_add_23_U36 ( .A(p11_C[54]), .B(
        p11_final_product2_25_), .ZN(p11_Partial_products_sum_add_23_n258) );
  NAND2_X1 p11_Partial_products_sum_add_23_U96 ( .A1(p11_C[35]), .A2(p11_S[36]), .ZN(p11_Partial_products_sum_add_23_n309) );
  NOR2_X1 p11_Partial_products_sum_add_23_U97 ( .A1(p11_C[35]), .A2(p11_S[36]), 
        .ZN(p11_Partial_products_sum_add_23_n308) );
  INV_X1 p9_Partial_products_sum_add_23_U40 ( .A(p9_C[53]), .ZN(
        p9_Partial_products_sum_add_23_n198) );
  INV_X1 p9_Partial_products_sum_add_23_U39 ( .A(p9_S[54]), .ZN(
        p9_Partial_products_sum_add_23_n197) );
  INV_X1 p9_Partial_products_sum_add_23_U48 ( .A(p9_C[51]), .ZN(
        p9_Partial_products_sum_add_23_n204) );
  INV_X1 p9_Partial_products_sum_add_23_U47 ( .A(p9_S[52]), .ZN(
        p9_Partial_products_sum_add_23_n203) );
  INV_X1 p9_Partial_products_sum_add_23_U56 ( .A(p9_C[49]), .ZN(
        p9_Partial_products_sum_add_23_n210) );
  INV_X1 p9_Partial_products_sum_add_23_U55 ( .A(p9_S[50]), .ZN(
        p9_Partial_products_sum_add_23_n209) );
  INV_X1 p9_Partial_products_sum_add_23_U64 ( .A(p9_C[47]), .ZN(
        p9_Partial_products_sum_add_23_n216) );
  INV_X1 p9_Partial_products_sum_add_23_U63 ( .A(p9_S[48]), .ZN(
        p9_Partial_products_sum_add_23_n215) );
  INV_X1 p9_Partial_products_sum_add_23_U72 ( .A(p9_C[45]), .ZN(
        p9_Partial_products_sum_add_23_n222) );
  INV_X1 p9_Partial_products_sum_add_23_U71 ( .A(p9_S[46]), .ZN(
        p9_Partial_products_sum_add_23_n221) );
  INV_X1 p9_Partial_products_sum_add_23_U80 ( .A(p9_C[43]), .ZN(
        p9_Partial_products_sum_add_23_n228) );
  INV_X1 p9_Partial_products_sum_add_23_U79 ( .A(p9_S[44]), .ZN(
        p9_Partial_products_sum_add_23_n227) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U82 ( .A(
        p9_Partial_products_sum_add_23_n231), .B(
        p9_Partial_products_sum_add_23_n230), .ZN(temp4[0]) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U109 ( .A(p9_S[43]), .B(p9_C[42]), 
        .ZN(p9_Partial_products_sum_add_23_n231) );
  AOI22_X1 p9_Partial_products_sum_add_23_U78 ( .A1(p9_S[44]), .A2(p9_C[43]), 
        .B1(p9_Partial_products_sum_add_23_n228), .B2(
        p9_Partial_products_sum_add_23_n227), .ZN(
        p9_Partial_products_sum_add_23_n229) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U76 ( .A(p9_S[45]), .B(p9_C[44]), 
        .ZN(p9_Partial_products_sum_add_23_n225) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U69 ( .A(
        p9_Partial_products_sum_add_23_n220), .B(
        p9_Partial_products_sum_add_23_n223), .ZN(temp4[3]) );
  AOI22_X1 p9_Partial_products_sum_add_23_U70 ( .A1(p9_S[46]), .A2(p9_C[45]), 
        .B1(p9_Partial_products_sum_add_23_n222), .B2(
        p9_Partial_products_sum_add_23_n221), .ZN(
        p9_Partial_products_sum_add_23_n223) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U68 ( .A(p9_S[47]), .B(p9_C[46]), 
        .ZN(p9_Partial_products_sum_add_23_n219) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U61 ( .A(
        p9_Partial_products_sum_add_23_n214), .B(
        p9_Partial_products_sum_add_23_n217), .ZN(temp4[5]) );
  AOI22_X1 p9_Partial_products_sum_add_23_U62 ( .A1(p9_S[48]), .A2(p9_C[47]), 
        .B1(p9_Partial_products_sum_add_23_n216), .B2(
        p9_Partial_products_sum_add_23_n215), .ZN(
        p9_Partial_products_sum_add_23_n217) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U60 ( .A(p9_S[49]), .B(p9_C[48]), 
        .ZN(p9_Partial_products_sum_add_23_n213) );
  AOI22_X1 p9_Partial_products_sum_add_23_U54 ( .A1(p9_S[50]), .A2(p9_C[49]), 
        .B1(p9_Partial_products_sum_add_23_n210), .B2(
        p9_Partial_products_sum_add_23_n209), .ZN(
        p9_Partial_products_sum_add_23_n211) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U52 ( .A(p9_S[51]), .B(p9_C[50]), 
        .ZN(p9_Partial_products_sum_add_23_n207) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U45 ( .A(
        p9_Partial_products_sum_add_23_n202), .B(
        p9_Partial_products_sum_add_23_n205), .ZN(temp4[9]) );
  AOI22_X1 p9_Partial_products_sum_add_23_U46 ( .A1(p9_S[52]), .A2(p9_C[51]), 
        .B1(p9_Partial_products_sum_add_23_n204), .B2(
        p9_Partial_products_sum_add_23_n203), .ZN(
        p9_Partial_products_sum_add_23_n205) );
  XNOR2_X1 p9_Partial_products_sum_add_23_U44 ( .A(p9_S[53]), .B(p9_C[52]), 
        .ZN(p9_Partial_products_sum_add_23_n201) );
  AOI22_X1 p9_Partial_products_sum_add_23_U38 ( .A1(p9_S[54]), .A2(p9_C[53]), 
        .B1(p9_Partial_products_sum_add_23_n198), .B2(
        p9_Partial_products_sum_add_23_n197), .ZN(
        p9_Partial_products_sum_add_23_n199) );
  OAI21_X1 p9_Partial_products_sum_add_23_U83 ( .B1(
        p9_Partial_products_sum_add_23_n232), .B2(
        p9_Partial_products_sum_add_23_n233), .A(
        p9_Partial_products_sum_add_23_n234), .ZN(
        p9_Partial_products_sum_add_23_n230) );
  NAND2_X1 p9_Partial_products_sum_add_23_U88 ( .A1(p9_C[39]), .A2(p9_S[40]), 
        .ZN(p9_Partial_products_sum_add_23_n238) );
  NOR2_X1 p9_Partial_products_sum_add_23_U89 ( .A1(p9_C[39]), .A2(p9_S[40]), 
        .ZN(p9_Partial_products_sum_add_23_n237) );
  NAND2_X1 p9_Partial_products_sum_add_23_U92 ( .A1(p9_C[37]), .A2(p9_S[38]), 
        .ZN(p9_Partial_products_sum_add_23_n242) );
  NOR2_X1 p9_Partial_products_sum_add_23_U93 ( .A1(p9_C[37]), .A2(p9_S[38]), 
        .ZN(p9_Partial_products_sum_add_23_n241) );
  NAND2_X1 p9_Partial_products_sum_add_23_U96 ( .A1(p9_C[35]), .A2(p9_S[36]), 
        .ZN(p9_Partial_products_sum_add_23_n246) );
  NOR2_X1 p9_Partial_products_sum_add_23_U97 ( .A1(p9_C[35]), .A2(p9_S[36]), 
        .ZN(p9_Partial_products_sum_add_23_n245) );
  NAND2_X1 p9_Partial_products_sum_add_23_U100 ( .A1(p9_S[34]), .A2(p9_C[33]), 
        .ZN(p9_Partial_products_sum_add_23_n250) );
  NOR2_X1 p9_Partial_products_sum_add_23_U101 ( .A1(p9_S[34]), .A2(p9_C[33]), 
        .ZN(p9_Partial_products_sum_add_23_n249) );
  NAND2_X1 p9_Partial_products_sum_add_23_U104 ( .A1(n3542), .A2(reg4_reg[3]), 
        .ZN(p9_Partial_products_sum_add_23_n253) );
  OAI21_X1 p9_Partial_products_sum_add_23_U105 ( .B1(n3542), .B2(reg4_reg[3]), 
        .A(p9_S[32]), .ZN(p9_Partial_products_sum_add_23_n252) );
  XOR2_X1 p9_Partial_products_sum_add_23_U110 ( .A(p9_final_product2_26_), .B(
        p9_final_product1_26), .Z(p9_Partial_products_sum_add_23_n193) );
  INV_X1 p8_Partial_products_sum_add_23_U40 ( .A(p8_C[53]), .ZN(
        p8_Partial_products_sum_add_23_n195) );
  INV_X1 p8_Partial_products_sum_add_23_U39 ( .A(p8_S[54]), .ZN(
        p8_Partial_products_sum_add_23_n194) );
  INV_X1 p8_Partial_products_sum_add_23_U56 ( .A(p8_C[49]), .ZN(
        p8_Partial_products_sum_add_23_n207) );
  INV_X1 p8_Partial_products_sum_add_23_U55 ( .A(p8_S[50]), .ZN(
        p8_Partial_products_sum_add_23_n206) );
  INV_X1 p8_Partial_products_sum_add_23_U64 ( .A(p8_C[47]), .ZN(
        p8_Partial_products_sum_add_23_n213) );
  INV_X1 p8_Partial_products_sum_add_23_U63 ( .A(p8_S[48]), .ZN(
        p8_Partial_products_sum_add_23_n212) );
  INV_X1 p8_Partial_products_sum_add_23_U72 ( .A(p8_C[45]), .ZN(
        p8_Partial_products_sum_add_23_n219) );
  INV_X1 p8_Partial_products_sum_add_23_U71 ( .A(p8_S[46]), .ZN(
        p8_Partial_products_sum_add_23_n218) );
  INV_X1 p8_Partial_products_sum_add_23_U80 ( .A(p8_C[43]), .ZN(
        p8_Partial_products_sum_add_23_n225) );
  INV_X1 p8_Partial_products_sum_add_23_U47 ( .A(p8_S[52]), .ZN(
        p8_Partial_products_sum_add_23_n200) );
  INV_X1 p8_Partial_products_sum_add_23_U48 ( .A(p8_C[51]), .ZN(
        p8_Partial_products_sum_add_23_n201) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U109 ( .A(p8_S[43]), .B(p8_C[42]), 
        .ZN(p8_Partial_products_sum_add_23_n228) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U76 ( .A(p8_S[45]), .B(p8_C[44]), 
        .ZN(p8_Partial_products_sum_add_23_n222) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U69 ( .A(
        p8_Partial_products_sum_add_23_n217), .B(
        p8_Partial_products_sum_add_23_n220), .ZN(temp3[3]) );
  AOI22_X1 p8_Partial_products_sum_add_23_U70 ( .A1(p8_S[46]), .A2(p8_C[45]), 
        .B1(p8_Partial_products_sum_add_23_n219), .B2(
        p8_Partial_products_sum_add_23_n218), .ZN(
        p8_Partial_products_sum_add_23_n220) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U68 ( .A(p8_S[47]), .B(p8_C[46]), 
        .ZN(p8_Partial_products_sum_add_23_n216) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U61 ( .A(
        p8_Partial_products_sum_add_23_n211), .B(
        p8_Partial_products_sum_add_23_n214), .ZN(temp3[5]) );
  AOI22_X1 p8_Partial_products_sum_add_23_U62 ( .A1(p8_S[48]), .A2(p8_C[47]), 
        .B1(p8_Partial_products_sum_add_23_n213), .B2(
        p8_Partial_products_sum_add_23_n212), .ZN(
        p8_Partial_products_sum_add_23_n214) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U60 ( .A(p8_S[49]), .B(p8_C[48]), 
        .ZN(p8_Partial_products_sum_add_23_n210) );
  AOI22_X1 p8_Partial_products_sum_add_23_U54 ( .A1(p8_S[50]), .A2(p8_C[49]), 
        .B1(p8_Partial_products_sum_add_23_n207), .B2(
        p8_Partial_products_sum_add_23_n206), .ZN(
        p8_Partial_products_sum_add_23_n208) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U52 ( .A(p8_S[51]), .B(p8_C[50]), 
        .ZN(p8_Partial_products_sum_add_23_n204) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U45 ( .A(
        p8_Partial_products_sum_add_23_n199), .B(
        p8_Partial_products_sum_add_23_n202), .ZN(temp3[9]) );
  AOI22_X1 p8_Partial_products_sum_add_23_U46 ( .A1(p8_S[52]), .A2(p8_C[51]), 
        .B1(p8_Partial_products_sum_add_23_n201), .B2(
        p8_Partial_products_sum_add_23_n200), .ZN(
        p8_Partial_products_sum_add_23_n202) );
  XNOR2_X1 p8_Partial_products_sum_add_23_U44 ( .A(p8_S[53]), .B(p8_C[52]), 
        .ZN(p8_Partial_products_sum_add_23_n198) );
  AOI22_X1 p8_Partial_products_sum_add_23_U38 ( .A1(p8_S[54]), .A2(p8_C[53]), 
        .B1(p8_Partial_products_sum_add_23_n195), .B2(
        p8_Partial_products_sum_add_23_n194), .ZN(
        p8_Partial_products_sum_add_23_n196) );
  AOI222_X1 p8_Partial_products_sum_add_23_U75 ( .A1(
        p8_Partial_products_sum_add_23_n223), .A2(
        p8_Partial_products_sum_add_23_n224), .B1(
        p8_Partial_products_sum_add_23_n223), .B2(
        p8_Partial_products_sum_add_23_n225), .C1(
        p8_Partial_products_sum_add_23_n224), .C2(
        p8_Partial_products_sum_add_23_n225), .ZN(
        p8_Partial_products_sum_add_23_n221) );
  NAND2_X1 p8_Partial_products_sum_add_23_U88 ( .A1(p8_C[39]), .A2(p8_S[40]), 
        .ZN(p8_Partial_products_sum_add_23_n235) );
  NOR2_X1 p8_Partial_products_sum_add_23_U89 ( .A1(p8_C[39]), .A2(p8_S[40]), 
        .ZN(p8_Partial_products_sum_add_23_n234) );
  NAND2_X1 p8_Partial_products_sum_add_23_U92 ( .A1(p8_C[37]), .A2(p8_S[38]), 
        .ZN(p8_Partial_products_sum_add_23_n239) );
  NOR2_X1 p8_Partial_products_sum_add_23_U93 ( .A1(p8_C[37]), .A2(p8_S[38]), 
        .ZN(p8_Partial_products_sum_add_23_n238) );
  NAND2_X1 p8_Partial_products_sum_add_23_U96 ( .A1(p8_C[35]), .A2(p8_S[36]), 
        .ZN(p8_Partial_products_sum_add_23_n243) );
  NOR2_X1 p8_Partial_products_sum_add_23_U97 ( .A1(p8_C[35]), .A2(p8_S[36]), 
        .ZN(p8_Partial_products_sum_add_23_n242) );
  NAND2_X1 p8_Partial_products_sum_add_23_U100 ( .A1(p8_S[34]), .A2(p8_C[33]), 
        .ZN(p8_Partial_products_sum_add_23_n247) );
  NAND2_X1 p8_Partial_products_sum_add_23_U104 ( .A1(n3511), .A2(reg3_reg[3]), 
        .ZN(p8_Partial_products_sum_add_23_n250) );
  OAI21_X1 p8_Partial_products_sum_add_23_U105 ( .B1(n3511), .B2(reg3_reg[3]), 
        .A(p8_S[32]), .ZN(p8_Partial_products_sum_add_23_n249) );
  XOR2_X1 p8_Partial_products_sum_add_23_U110 ( .A(p8_final_product2_26_), .B(
        p8_final_product1_26), .Z(p8_Partial_products_sum_add_23_n190) );
  INV_X1 p7_Partial_products_sum_add_23_U40 ( .A(p7_C[53]), .ZN(
        p7_Partial_products_sum_add_23_n195) );
  INV_X1 p7_Partial_products_sum_add_23_U39 ( .A(p7_S[54]), .ZN(
        p7_Partial_products_sum_add_23_n194) );
  INV_X1 p7_Partial_products_sum_add_23_U48 ( .A(p7_C[51]), .ZN(
        p7_Partial_products_sum_add_23_n201) );
  INV_X1 p7_Partial_products_sum_add_23_U47 ( .A(p7_S[52]), .ZN(
        p7_Partial_products_sum_add_23_n200) );
  INV_X1 p7_Partial_products_sum_add_23_U56 ( .A(p7_C[49]), .ZN(
        p7_Partial_products_sum_add_23_n207) );
  INV_X1 p7_Partial_products_sum_add_23_U55 ( .A(p7_S[50]), .ZN(
        p7_Partial_products_sum_add_23_n206) );
  INV_X1 p7_Partial_products_sum_add_23_U64 ( .A(p7_C[47]), .ZN(
        p7_Partial_products_sum_add_23_n213) );
  INV_X1 p7_Partial_products_sum_add_23_U63 ( .A(p7_S[48]), .ZN(
        p7_Partial_products_sum_add_23_n212) );
  INV_X1 p7_Partial_products_sum_add_23_U72 ( .A(p7_C[45]), .ZN(
        p7_Partial_products_sum_add_23_n219) );
  INV_X1 p7_Partial_products_sum_add_23_U71 ( .A(p7_S[46]), .ZN(
        p7_Partial_products_sum_add_23_n218) );
  INV_X1 p7_Partial_products_sum_add_23_U80 ( .A(p7_C[43]), .ZN(
        p7_Partial_products_sum_add_23_n225) );
  INV_X1 p7_Partial_products_sum_add_23_U79 ( .A(p7_S[44]), .ZN(
        p7_Partial_products_sum_add_23_n224) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U82 ( .A(
        p7_Partial_products_sum_add_23_n228), .B(
        p7_Partial_products_sum_add_23_n227), .ZN(temp2[0]) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U109 ( .A(p7_S[43]), .B(p7_C[42]), 
        .ZN(p7_Partial_products_sum_add_23_n228) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U77 ( .A(
        p7_Partial_products_sum_add_23_n223), .B(
        p7_Partial_products_sum_add_23_n226), .ZN(temp2[1]) );
  AOI22_X1 p7_Partial_products_sum_add_23_U78 ( .A1(p7_S[44]), .A2(p7_C[43]), 
        .B1(p7_Partial_products_sum_add_23_n225), .B2(
        p7_Partial_products_sum_add_23_n224), .ZN(
        p7_Partial_products_sum_add_23_n226) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U76 ( .A(p7_S[45]), .B(p7_C[44]), 
        .ZN(p7_Partial_products_sum_add_23_n222) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U69 ( .A(
        p7_Partial_products_sum_add_23_n217), .B(
        p7_Partial_products_sum_add_23_n220), .ZN(temp2[3]) );
  AOI22_X1 p7_Partial_products_sum_add_23_U70 ( .A1(p7_S[46]), .A2(p7_C[45]), 
        .B1(p7_Partial_products_sum_add_23_n219), .B2(
        p7_Partial_products_sum_add_23_n218), .ZN(
        p7_Partial_products_sum_add_23_n220) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U68 ( .A(p7_S[47]), .B(p7_C[46]), 
        .ZN(p7_Partial_products_sum_add_23_n216) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U61 ( .A(
        p7_Partial_products_sum_add_23_n211), .B(
        p7_Partial_products_sum_add_23_n214), .ZN(temp2[5]) );
  AOI22_X1 p7_Partial_products_sum_add_23_U62 ( .A1(p7_S[48]), .A2(p7_C[47]), 
        .B1(p7_Partial_products_sum_add_23_n213), .B2(
        p7_Partial_products_sum_add_23_n212), .ZN(
        p7_Partial_products_sum_add_23_n214) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U60 ( .A(p7_S[49]), .B(p7_C[48]), 
        .ZN(p7_Partial_products_sum_add_23_n210) );
  AOI22_X1 p7_Partial_products_sum_add_23_U54 ( .A1(p7_S[50]), .A2(p7_C[49]), 
        .B1(p7_Partial_products_sum_add_23_n207), .B2(
        p7_Partial_products_sum_add_23_n206), .ZN(
        p7_Partial_products_sum_add_23_n208) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U52 ( .A(p7_S[51]), .B(p7_C[50]), 
        .ZN(p7_Partial_products_sum_add_23_n204) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U45 ( .A(
        p7_Partial_products_sum_add_23_n199), .B(
        p7_Partial_products_sum_add_23_n202), .ZN(temp2[9]) );
  AOI22_X1 p7_Partial_products_sum_add_23_U46 ( .A1(p7_S[52]), .A2(p7_C[51]), 
        .B1(p7_Partial_products_sum_add_23_n201), .B2(
        p7_Partial_products_sum_add_23_n200), .ZN(
        p7_Partial_products_sum_add_23_n202) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U44 ( .A(p7_S[53]), .B(p7_C[52]), 
        .ZN(p7_Partial_products_sum_add_23_n198) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U37 ( .A(
        p7_Partial_products_sum_add_23_n193), .B(
        p7_Partial_products_sum_add_23_n196), .ZN(temp2[11]) );
  AOI22_X1 p7_Partial_products_sum_add_23_U38 ( .A1(p7_S[54]), .A2(p7_C[53]), 
        .B1(p7_Partial_products_sum_add_23_n195), .B2(
        p7_Partial_products_sum_add_23_n194), .ZN(
        p7_Partial_products_sum_add_23_n196) );
  XNOR2_X1 p7_Partial_products_sum_add_23_U36 ( .A(p7_C[54]), .B(
        p7_final_product2_25_), .ZN(p7_Partial_products_sum_add_23_n192) );
  NAND2_X1 p7_Partial_products_sum_add_23_U88 ( .A1(p7_C[39]), .A2(p7_S[40]), 
        .ZN(p7_Partial_products_sum_add_23_n235) );
  NOR2_X1 p7_Partial_products_sum_add_23_U89 ( .A1(p7_C[39]), .A2(p7_S[40]), 
        .ZN(p7_Partial_products_sum_add_23_n234) );
  NAND2_X1 p7_Partial_products_sum_add_23_U92 ( .A1(p7_C[37]), .A2(p7_S[38]), 
        .ZN(p7_Partial_products_sum_add_23_n239) );
  NOR2_X1 p7_Partial_products_sum_add_23_U93 ( .A1(p7_C[37]), .A2(p7_S[38]), 
        .ZN(p7_Partial_products_sum_add_23_n238) );
  NAND2_X1 p7_Partial_products_sum_add_23_U96 ( .A1(p7_C[35]), .A2(p7_S[36]), 
        .ZN(p7_Partial_products_sum_add_23_n243) );
  NOR2_X1 p7_Partial_products_sum_add_23_U97 ( .A1(p7_C[35]), .A2(p7_S[36]), 
        .ZN(p7_Partial_products_sum_add_23_n242) );
  NAND2_X1 p7_Partial_products_sum_add_23_U104 ( .A1(n3499), .A2(reg2_reg[3]), 
        .ZN(p7_Partial_products_sum_add_23_n250) );
  OAI21_X1 p7_Partial_products_sum_add_23_U105 ( .B1(n3499), .B2(reg2_reg[3]), 
        .A(p7_S[32]), .ZN(p7_Partial_products_sum_add_23_n249) );
  XOR2_X1 p7_Partial_products_sum_add_23_U110 ( .A(p7_final_product2_26_), .B(
        p7_final_product1_26), .Z(p7_Partial_products_sum_add_23_n190) );
  DFFS_X1 REGISTER4_q_reg_10_ ( .D(n3272), .CK(CLK), .SN(RST_n), .QN(
        reg4_reg[10]) );
  DFFR_X1 REG11_q_reg_12_ ( .D(REG11_n49), .CK(CLK), .RN(RST_n), .Q(reg2[12]), 
        .QN(n3690) );
  DFFR_X1 REG11_q_reg_11_ ( .D(REG11_n50), .CK(CLK), .RN(RST_n), .Q(reg2[11]), 
        .QN(n3686) );
  DFFR_X1 REG11_q_reg_8_ ( .D(REG11_n53), .CK(CLK), .RN(RST_n), .Q(reg2[8]), 
        .QN(n3683) );
  DFFR_X1 REGISTER4_q_reg_1_ ( .D(REGISTER4_n60), .CK(CLK), .RN(RST_n), .Q(
        reg4_reg[1]), .QN(n3701) );
  DFFR_X1 REGISTER3_q_reg_1_ ( .D(REGISTER3_n60), .CK(CLK), .RN(RST_n), .Q(
        reg3_reg[1]), .QN(n3700) );
  DFFR_X1 REGISTER2_q_reg_1_ ( .D(REGISTER2_n60), .CK(CLK), .RN(RST_n), .Q(
        reg2_reg[1]), .QN(n3716) );
  AOI221_X1 U3434 ( .B1(n2497), .B2(reg2[1]), .C1(n2498), .C2(n3684), .A(n2752), .ZN(n2407) );
  AOI221_X1 U3435 ( .B1(n2047), .B2(B0[3]), .C1(n2048), .C2(n2115), .A(n2273), 
        .ZN(n2253) );
  AOI221_X1 U3436 ( .B1(n2047), .B2(B0[2]), .C1(n2048), .C2(n2133), .A(n2282), 
        .ZN(n2262) );
  AOI221_X1 U3437 ( .B1(n2497), .B2(reg2[3]), .C1(n2498), .C2(n3669), .A(n2725), .ZN(n2705) );
  AOI222_X1 U3438 ( .A1(n2401), .A2(n2402), .B1(n2401), .B2(n2399), .C1(n2402), 
        .C2(n2399), .ZN(p11_C[39]) );
  AOI221_X1 U3439 ( .B1(n2947), .B2(reg4[12]), .C1(n2948), .C2(n3679), .A(
        n2970), .ZN(n2949) );
  AOI221_X1 U3440 ( .B1(n2947), .B2(reg4[11]), .C1(n2948), .C2(n3671), .A(
        n2986), .ZN(n2971) );
  AOI221_X1 U3441 ( .B1(n2497), .B2(reg2[9]), .C1(n2498), .C2(n3691), .A(n2598), .ZN(n2554) );
  AOI221_X1 U3442 ( .B1(n2497), .B2(reg2[8]), .C1(n2498), .C2(n3683), .A(n2627), .ZN(n2626) );
  AOI221_X1 U3443 ( .B1(n2497), .B2(reg2[7]), .C1(n2498), .C2(n3688), .A(n2639), .ZN(n2612) );
  INV_X1 U3444 ( .A(B0[10]), .ZN(n1991) );
  AOI222_X1 U3445 ( .A1(n1008), .A2(n1009), .B1(n1008), .B2(n1006), .C1(n1009), 
        .C2(n1006), .ZN(p8_C[50]) );
  AOI222_X1 U3446 ( .A1(n1040), .A2(n1041), .B1(n1040), .B2(n1038), .C1(n1041), 
        .C2(n1038), .ZN(p8_C[42]) );
  AOI22_X1 U3447 ( .A1(n1997), .A2(B0[9]), .B1(n1996), .B2(n2003), .ZN(n3339)
         );
  AND2_X1 U3448 ( .A1(n2006), .A2(B0[10]), .ZN(n3340) );
  AOI211_X1 U3449 ( .C1(n1991), .C2(n2007), .A(n3339), .B(n3340), .ZN(n2052)
         );
  AOI22_X1 U3450 ( .A1(n2922), .A2(reg4[9]), .B1(n2921), .B2(n3681), .ZN(n3341) );
  AND2_X1 U3451 ( .A1(n2947), .A2(reg4[10]), .ZN(n3342) );
  AOI211_X1 U3452 ( .C1(n3682), .C2(n2948), .A(n3341), .B(n3342), .ZN(n2979)
         );
  AND2_X1 U3453 ( .A1(n3687), .A2(n2498), .ZN(n3343) );
  AOI22_X1 U3454 ( .A1(reg2[5]), .A2(n3662), .B1(n3677), .B2(n2471), .ZN(n3344) );
  AOI211_X1 U3455 ( .C1(reg2[6]), .C2(n2497), .A(n3343), .B(n3344), .ZN(n2644)
         );
  OAI21_X1 U3456 ( .B1(A1[2]), .B2(A1[1]), .A(A1[3]), .ZN(n3345) );
  AOI21_X2 U3457 ( .B1(A1[2]), .B2(A1[1]), .A(n3345), .ZN(n2602) );
  OAI22_X1 U3458 ( .A1(n1889), .A2(n1888), .B1(n1887), .B2(B0[0]), .ZN(n3346)
         );
  INV_X1 U3459 ( .A(n3346), .ZN(n3347) );
  AOI222_X1 U3460 ( .A1(B0[1]), .A2(n1884), .B1(n1888), .B2(n3777), .C1(n1885), 
        .C2(n1886), .ZN(n3348) );
  INV_X1 U3461 ( .A(reg1_reg[1]), .ZN(n3349) );
  AOI211_X1 U3462 ( .C1(n1882), .C2(n3347), .A(n3348), .B(n3349), .ZN(n3654)
         );
  INV_X1 U3463 ( .A(A2[3]), .ZN(n3350) );
  XNOR2_X1 U3464 ( .A(n2878), .B(n2877), .ZN(n3351) );
  AOI22_X1 U3465 ( .A1(n2784), .A2(reg4[1]), .B1(n3666), .B2(n2785), .ZN(n3352) );
  OAI21_X1 U3466 ( .B1(reg4[0]), .B2(n2782), .A(n3352), .ZN(n3353) );
  NAND3_X1 U3467 ( .A1(\p10/final_product1[0] ), .A2(A2[1]), .A3(n3353), .ZN(
        n3354) );
  AOI222_X1 U3468 ( .A1(n3350), .A2(n3351), .B1(n3350), .B2(n3354), .C1(n3351), 
        .C2(n3354), .ZN(p10_Partial_products_sum_add_23_n340) );
  AND2_X1 U3469 ( .A1(n2041), .A2(n2048), .ZN(n3355) );
  AOI22_X1 U3470 ( .A1(B0[5]), .A2(n2022), .B1(n2063), .B2(n2021), .ZN(n3356)
         );
  AOI211_X1 U3471 ( .C1(n2047), .C2(B0[6]), .A(n3355), .B(n3356), .ZN(n2191)
         );
  NAND2_X1 U3472 ( .A1(n1821), .A2(n1820), .ZN(n3357) );
  XOR2_X1 U3473 ( .A(n1806), .B(n3357), .Z(n1808) );
  AOI22_X1 U3474 ( .A1(n2922), .A2(reg4[8]), .B1(n2921), .B2(n3667), .ZN(n3358) );
  AND2_X1 U3475 ( .A1(n2947), .A2(reg4[9]), .ZN(n3359) );
  AOI211_X1 U3476 ( .C1(n3681), .C2(n2948), .A(n3358), .B(n3359), .ZN(n3003)
         );
  AOI22_X1 U3477 ( .A1(n3826), .A2(reg2[7]), .B1(n2517), .B2(n3688), .ZN(n3360) );
  AND2_X1 U3478 ( .A1(n2531), .A2(reg2[8]), .ZN(n3361) );
  AOI211_X1 U3479 ( .C1(n3683), .C2(n2532), .A(n3360), .B(n3361), .ZN(n2635)
         );
  AND2_X1 U3480 ( .A1(n3685), .A2(n2498), .ZN(n3362) );
  AOI22_X1 U3481 ( .A1(reg2[3]), .A2(n3662), .B1(n3669), .B2(n2471), .ZN(n3363) );
  AOI211_X1 U3482 ( .C1(reg2[4]), .C2(n2497), .A(n3362), .B(n3363), .ZN(n2685)
         );
  AOI22_X1 U3483 ( .A1(n3689), .A2(n2532), .B1(reg2[0]), .B2(n2531), .ZN(n3364) );
  AND2_X1 U3484 ( .A1(n2517), .A2(n3364), .ZN(n2424) );
  NAND2_X1 U3485 ( .A1(n1977), .A2(n1978), .ZN(n3365) );
  OAI221_X1 U3486 ( .B1(n3654), .B2(reg1_reg[3]), .C1(n1977), .C2(n1978), .A(
        n3365), .ZN(p6_Partial_products_sum_add_23_n232) );
  XOR2_X1 U3487 ( .A(n1521), .B(n1522), .Z(n3366) );
  OR2_X1 U3488 ( .A1(n1525), .A2(n1526), .ZN(n3367) );
  AOI222_X1 U3489 ( .A1(p7_Partial_products_sum_add_23_n248), .A2(p7_C[32]), 
        .B1(p7_Partial_products_sum_add_23_n248), .B2(p7_S[33]), .C1(p7_C[32]), 
        .C2(p7_S[33]), .ZN(n3368) );
  AOI222_X1 U3490 ( .A1(n3366), .A2(n3367), .B1(n3366), .B2(n3368), .C1(n3367), 
        .C2(n3368), .ZN(p7_Partial_products_sum_add_23_n244) );
  OAI21_X1 U3491 ( .B1(p8_Partial_products_sum_add_23_n240), .B2(p8_C[36]), 
        .A(p8_S[37]), .ZN(n3369) );
  AND2_X1 U3492 ( .A1(n3369), .A2(n3502), .ZN(
        p8_Partial_products_sum_add_23_n237) );
  AOI22_X1 U3493 ( .A1(n2922), .A2(reg4[0]), .B1(n2921), .B2(n3670), .ZN(n3370) );
  AND2_X1 U3494 ( .A1(n2947), .A2(reg4[1]), .ZN(n3371) );
  AOI211_X1 U3495 ( .C1(n3666), .C2(n2948), .A(n3370), .B(n3371), .ZN(n2857)
         );
  NAND2_X1 U3496 ( .A1(n2270), .A2(n2271), .ZN(n3372) );
  XOR2_X1 U3497 ( .A(n2256), .B(n3372), .Z(n2258) );
  AOI22_X1 U3498 ( .A1(n2022), .A2(B0[3]), .B1(n2021), .B2(n2115), .ZN(n3373)
         );
  AND2_X1 U3499 ( .A1(n2047), .A2(B0[4]), .ZN(n3374) );
  AOI211_X1 U3500 ( .C1(n2075), .C2(n2048), .A(n3373), .B(n3374), .ZN(n2233)
         );
  NAND2_X1 U3501 ( .A1(n1801), .A2(n1800), .ZN(n3375) );
  XOR2_X1 U3502 ( .A(n1775), .B(n3375), .Z(n1777) );
  OAI21_X1 U3503 ( .B1(p7_Partial_products_sum_add_23_n236), .B2(p7_C[38]), 
        .A(p7_S[39]), .ZN(n3376) );
  AND2_X1 U3504 ( .A1(n3376), .A2(n3489), .ZN(
        p7_Partial_products_sum_add_23_n233) );
  XOR2_X1 U3505 ( .A(n1324), .B(reg3_reg[11]), .Z(n1046) );
  AOI22_X1 U3506 ( .A1(n1169), .A2(B2[6]), .B1(n1168), .B2(n1142), .ZN(n3377)
         );
  AND2_X1 U3507 ( .A1(n1182), .A2(B2[7]), .ZN(n3378) );
  AOI211_X1 U3508 ( .C1(n1118), .C2(n1183), .A(n3377), .B(n3378), .ZN(n1320)
         );
  AOI22_X1 U3509 ( .A1(n3048), .A2(n3682), .B1(n3047), .B2(reg4[10]), .ZN(
        n3379) );
  OR2_X1 U3510 ( .A1(n3836), .A2(reg4[9]), .ZN(n3380) );
  OAI211_X1 U3511 ( .C1(n3009), .C2(n3681), .A(n3379), .B(n3380), .ZN(n3381)
         );
  XNOR2_X1 U3512 ( .A(n3080), .B(n3381), .ZN(n3082) );
  XOR2_X1 U3513 ( .A(n3122), .B(A2[11]), .Z(n2845) );
  INV_X1 U3514 ( .A(A1[2]), .ZN(n3382) );
  INV_X1 U3515 ( .A(A1[1]), .ZN(n3383) );
  AOI221_X4 U3516 ( .B1(A1[2]), .B2(A1[1]), .C1(n3382), .C2(n3383), .A(A1[3]), 
        .ZN(n2601) );
  INV_X1 U3517 ( .A(n2614), .ZN(n3384) );
  AOI22_X1 U3518 ( .A1(n2614), .A2(n2613), .B1(n2612), .B2(n3384), .ZN(n2583)
         );
  INV_X1 U3519 ( .A(n1432), .ZN(n3385) );
  AOI222_X1 U3520 ( .A1(n3385), .A2(n1438), .B1(n1436), .B2(n1435), .C1(B1[1]), 
        .C2(n1434), .ZN(n3386) );
  INV_X1 U3521 ( .A(n3386), .ZN(p7_final_product1[1]) );
  AOI22_X1 U3522 ( .A1(n3670), .A2(n2985), .B1(reg4[0]), .B2(n2984), .ZN(n3387) );
  AND2_X1 U3523 ( .A1(n2967), .A2(n3387), .ZN(n2874) );
  XOR2_X1 U3524 ( .A(n1963), .B(n1964), .Z(n1967) );
  OAI21_X1 U3525 ( .B1(p8_S[35]), .B2(p8_C[34]), .A(
        p8_Partial_products_sum_add_23_n244), .ZN(n3388) );
  AND2_X1 U3526 ( .A1(n3388), .A2(n3501), .ZN(
        p8_Partial_products_sum_add_23_n241) );
  OAI21_X1 U3527 ( .B1(p7_Partial_products_sum_add_23_n240), .B2(p7_C[36]), 
        .A(p7_S[37]), .ZN(n3389) );
  AND2_X1 U3528 ( .A1(n3389), .A2(n3487), .ZN(
        p7_Partial_products_sum_add_23_n237) );
  OAI21_X1 U3529 ( .B1(p9_Partial_products_sum_add_23_n243), .B2(p9_C[36]), 
        .A(p9_S[37]), .ZN(n3390) );
  AND2_X1 U3530 ( .A1(n3390), .A2(n3524), .ZN(
        p9_Partial_products_sum_add_23_n240) );
  XOR2_X1 U3531 ( .A(n3721), .B(n1361), .Z(n1055) );
  AOI22_X1 U3532 ( .A1(B0[10]), .A2(n2148), .B1(n1991), .B2(n2149), .ZN(n3391)
         );
  OAI211_X1 U3533 ( .C1(B0[9]), .C2(n2111), .A(n3832), .B(n3391), .ZN(n3392)
         );
  XNOR2_X1 U3534 ( .A(n2180), .B(n3392), .ZN(n2182) );
  XOR2_X1 U3535 ( .A(reg1_reg[11]), .B(n2224), .Z(n1945) );
  NAND2_X1 U3536 ( .A1(n3148), .A2(n3149), .ZN(n3393) );
  XOR2_X1 U3537 ( .A(n3123), .B(n3393), .Z(n3125) );
  AOI22_X1 U3538 ( .A1(n3662), .A2(reg2[11]), .B1(n2471), .B2(n3686), .ZN(
        n3394) );
  AND2_X1 U3539 ( .A1(n2497), .A2(reg2[12]), .ZN(n3395) );
  AOI211_X1 U3540 ( .C1(n3690), .C2(n2498), .A(n3394), .B(n3395), .ZN(n2499)
         );
  XOR2_X1 U3541 ( .A(n2130), .B(n2123), .Z(n3396) );
  XNOR2_X1 U3542 ( .A(n2124), .B(n3396), .ZN(n2131) );
  XOR2_X1 U3543 ( .A(reg2_reg[11]), .B(n1774), .Z(n1495) );
  XOR2_X1 U3544 ( .A(n1301), .B(n1302), .Z(n1044) );
  AOI222_X1 U3545 ( .A1(n1320), .A2(n1318), .B1(n1320), .B2(n1319), .C1(n1318), 
        .C2(n1319), .ZN(n3397) );
  XOR2_X1 U3546 ( .A(n1298), .B(n3397), .Z(n1299) );
  XOR2_X1 U3547 ( .A(n843), .B(n844), .Z(n848) );
  NAND2_X1 U3548 ( .A1(p10_S[39]), .A2(p10_C[38]), .ZN(n3398) );
  NAND3_X1 U3549 ( .A1(n3398), .A2(n3579), .A3(n3578), .ZN(n3399) );
  OAI21_X1 U3550 ( .B1(n3399), .B2(p10_S[40]), .A(p10_C[39]), .ZN(n3400) );
  NAND2_X1 U3551 ( .A1(n3399), .A2(p10_S[40]), .ZN(n3401) );
  NAND2_X1 U3552 ( .A1(n3400), .A2(n3401), .ZN(
        p10_Partial_products_sum_add_23_n322) );
  AOI22_X1 U3553 ( .A1(n2922), .A2(reg4[4]), .B1(n2921), .B2(n3668), .ZN(n3402) );
  AND2_X1 U3554 ( .A1(n2947), .A2(reg4[5]), .ZN(n3403) );
  AOI211_X1 U3555 ( .C1(n3664), .C2(n2948), .A(n3402), .B(n3403), .ZN(n3102)
         );
  OAI21_X1 U3556 ( .B1(p11_Partial_products_sum_add_23_n260), .B2(
        p11_Partial_products_sum_add_23_n261), .A(
        p11_Partial_products_sum_add_23_n259), .ZN(n3564) );
  OAI22_X1 U3557 ( .A1(reg2[7]), .A2(n2561), .B1(reg2[9]), .B2(n2332), .ZN(
        n3404) );
  AOI22_X1 U3558 ( .A1(n3693), .A2(n2335), .B1(reg2[10]), .B2(n2334), .ZN(
        n3405) );
  AOI22_X1 U3559 ( .A1(reg2[8]), .A2(n2601), .B1(n3683), .B2(n2602), .ZN(n3406) );
  OAI211_X1 U3560 ( .C1(n3688), .C2(n2562), .A(n3405), .B(n3406), .ZN(n3407)
         );
  NOR2_X1 U3561 ( .A1(n3404), .A2(n3407), .ZN(n3408) );
  AOI21_X1 U3562 ( .B1(n2685), .B2(n2686), .A(n3408), .ZN(n3409) );
  XNOR2_X1 U3563 ( .A(n3409), .B(n2655), .ZN(n2657) );
  INV_X1 U3564 ( .A(n3761), .ZN(n3410) );
  NAND2_X1 U3565 ( .A1(B2[13]), .A2(n977), .ZN(n3411) );
  OAI22_X1 U3566 ( .A1(B2[13]), .A2(n3410), .B1(n979), .B2(n3411), .ZN(
        p8_final_product1_26) );
  OAI21_X1 U3567 ( .B1(p9_final_product2_25_), .B2(n3527), .A(p9_C[54]), .ZN(
        n3412) );
  AND2_X1 U3568 ( .A1(n3412), .A2(n3526), .ZN(
        p9_Partial_products_sum_add_23_n192) );
  XOR2_X1 U3569 ( .A(n2383), .B(n2385), .Z(n3413) );
  XNOR2_X1 U3570 ( .A(n2386), .B(n3413), .ZN(p11_S[43]) );
  INV_X1 U3571 ( .A(mul3_reg[12]), .ZN(n3414) );
  AOI222_X1 U3572 ( .A1(p8_Partial_products_sum_add_23_n195), .A2(
        p8_Partial_products_sum_add_23_n194), .B1(
        p8_Partial_products_sum_add_23_n195), .B2(
        p8_Partial_products_sum_add_23_n193), .C1(
        p8_Partial_products_sum_add_23_n194), .C2(
        p8_Partial_products_sum_add_23_n193), .ZN(n3415) );
  XOR2_X1 U3573 ( .A(p8_C[54]), .B(p8_final_product2_25_), .Z(n3416) );
  XNOR2_X1 U3574 ( .A(n3415), .B(n3416), .ZN(n3417) );
  INV_X1 U3575 ( .A(n3847), .ZN(n3418) );
  AOI22_X1 U3576 ( .A1(n3847), .A2(n3414), .B1(n3417), .B2(n3418), .ZN(
        REG3_1_n50) );
  OAI22_X1 U3577 ( .A1(n990), .A2(n989), .B1(n988), .B2(B2[0]), .ZN(n3419) );
  INV_X1 U3578 ( .A(n3419), .ZN(n3420) );
  AOI222_X1 U3579 ( .A1(B2[1]), .A2(n985), .B1(n989), .B2(n3816), .C1(n986), 
        .C2(n987), .ZN(n3421) );
  INV_X1 U3580 ( .A(reg3_reg[1]), .ZN(n3422) );
  AOI211_X1 U3581 ( .C1(n983), .C2(n3420), .A(n3421), .B(n3422), .ZN(n3511) );
  OAI22_X1 U3582 ( .A1(n540), .A2(n539), .B1(n538), .B2(B3[0]), .ZN(n3423) );
  INV_X1 U3583 ( .A(n3423), .ZN(n3424) );
  AOI222_X1 U3584 ( .A1(B3[1]), .A2(n535), .B1(n539), .B2(n3812), .C1(n536), 
        .C2(n537), .ZN(n3425) );
  INV_X1 U3585 ( .A(reg4_reg[1]), .ZN(n3426) );
  AOI211_X1 U3586 ( .C1(n533), .C2(n3424), .A(n3425), .B(n3426), .ZN(n3542) );
  OAI21_X1 U3587 ( .B1(p7_S[35]), .B2(p7_C[34]), .A(
        p7_Partial_products_sum_add_23_n244), .ZN(n3427) );
  AND2_X1 U3588 ( .A1(n3427), .A2(n3486), .ZN(
        p7_Partial_products_sum_add_23_n241) );
  OAI21_X1 U3589 ( .B1(p9_S[35]), .B2(p9_C[34]), .A(
        p9_Partial_products_sum_add_23_n247), .ZN(n3428) );
  AND2_X1 U3590 ( .A1(n3428), .A2(n3523), .ZN(
        p9_Partial_products_sum_add_23_n244) );
  AOI222_X1 U3591 ( .A1(B0[8]), .A2(n1884), .B1(n1885), .B2(n2005), .C1(n3777), 
        .C2(n2017), .ZN(n3429) );
  INV_X1 U3592 ( .A(n3429), .ZN(n2270) );
  AOI22_X1 U3593 ( .A1(n2048), .A2(n1888), .B1(n2047), .B2(B0[0]), .ZN(n3430)
         );
  AND2_X1 U3594 ( .A1(n2021), .A2(n3430), .ZN(n2293) );
  XOR2_X1 U3595 ( .A(n3719), .B(n1811), .Z(n1504) );
  XOR2_X1 U3596 ( .A(n3720), .B(n912), .Z(n605) );
  NAND2_X1 U3597 ( .A1(n2702), .A2(n2703), .ZN(n3431) );
  XOR2_X1 U3598 ( .A(n2677), .B(n3431), .Z(n2679) );
  AND2_X1 U3599 ( .A1(n1142), .A2(n1149), .ZN(n3432) );
  AOI22_X1 U3600 ( .A1(B2[5]), .A2(n1123), .B1(n1164), .B2(n1122), .ZN(n3433)
         );
  AOI211_X1 U3601 ( .C1(B2[6]), .C2(n1148), .A(n3432), .B(n3433), .ZN(n1292)
         );
  AOI22_X1 U3602 ( .A1(n1980), .A2(B0[9]), .B1(n1979), .B2(n2003), .ZN(n3434)
         );
  AND2_X1 U3603 ( .A1(n1988), .A2(B0[10]), .ZN(n3435) );
  AOI211_X1 U3604 ( .C1(n1991), .C2(n1989), .A(n3434), .B(n3435), .ZN(n2013)
         );
  XOR2_X1 U3605 ( .A(n2192), .B(n2193), .Z(n2197) );
  XOR2_X1 U3606 ( .A(n1750), .B(n1751), .Z(n1493) );
  XOR2_X1 U3607 ( .A(n3758), .B(n1745), .Z(n1489) );
  XNOR2_X1 U3608 ( .A(n1297), .B(n1307), .ZN(n1296) );
  XOR2_X1 U3609 ( .A(n875), .B(reg4_reg[11]), .Z(n596) );
  OAI21_X1 U3610 ( .B1(n3118), .B2(n3117), .A(n3116), .ZN(n3436) );
  NAND2_X1 U3611 ( .A1(n3436), .A2(n3817), .ZN(n3437) );
  XNOR2_X1 U3612 ( .A(n3096), .B(n3437), .ZN(n3097) );
  AOI222_X1 U3613 ( .A1(n2672), .A2(n2670), .B1(n2672), .B2(n2671), .C1(n2670), 
        .C2(n2671), .ZN(n3438) );
  XOR2_X1 U3614 ( .A(n2650), .B(n3438), .Z(n2651) );
  AOI22_X1 U3615 ( .A1(n3662), .A2(reg2[4]), .B1(n2471), .B2(n3685), .ZN(n3439) );
  AND2_X1 U3616 ( .A1(n2497), .A2(reg2[5]), .ZN(n3440) );
  AOI211_X1 U3617 ( .C1(n3677), .C2(n2498), .A(n3439), .B(n3440), .ZN(n2656)
         );
  OAI21_X1 U3618 ( .B1(p8_Partial_products_sum_add_23_n232), .B2(p8_C[40]), 
        .A(p8_S[41]), .ZN(n3441) );
  AND2_X1 U3619 ( .A1(n3441), .A2(n3503), .ZN(
        p8_Partial_products_sum_add_23_n229) );
  XOR2_X1 U3620 ( .A(n3773), .B(n846), .Z(n590) );
  MUX2_X1 U3621 ( .A(n3052), .B(n3053), .S(n3054), .Z(n2829) );
  INV_X1 U3622 ( .A(n1900), .ZN(n3442) );
  AOI222_X1 U3623 ( .A1(n1992), .A2(n1898), .B1(n1992), .B2(n3442), .C1(n1898), 
        .C2(n3442), .ZN(p6_C[52]) );
  NAND3_X1 U3624 ( .A1(n3639), .A2(n3637), .A3(n3638), .ZN(n3443) );
  OAI21_X1 U3625 ( .B1(n3443), .B2(p6_S[42]), .A(p6_C[41]), .ZN(n3444) );
  NAND2_X1 U3626 ( .A1(n3443), .A2(p6_S[42]), .ZN(n3445) );
  NAND2_X1 U3627 ( .A1(n3444), .A2(n3445), .ZN(
        p6_Partial_products_sum_add_23_n210) );
  OAI21_X1 U3628 ( .B1(p8_C[54]), .B2(n3504), .A(p8_final_product2_25_), .ZN(
        n3446) );
  AND2_X1 U3629 ( .A1(n3446), .A2(n3505), .ZN(
        p8_Partial_products_sum_add_23_n189) );
  OAI21_X1 U3630 ( .B1(p8_Partial_products_sum_add_23_n205), .B2(
        p8_Partial_products_sum_add_23_n207), .A(
        p8_Partial_products_sum_add_23_n206), .ZN(n3447) );
  AND2_X1 U3631 ( .A1(n3447), .A2(n3515), .ZN(
        p8_Partial_products_sum_add_23_n203) );
  NAND2_X1 U3632 ( .A1(fb_0_), .A2(xin[0]), .ZN(n3448) );
  OAI211_X1 U3633 ( .C1(fb_0_), .C2(xin[0]), .A(VIN), .B(n3448), .ZN(n3309) );
  OAI21_X1 U3634 ( .B1(p10_Partial_products_sum_add_23_n280), .B2(p10_C[53]), 
        .A(p10_S[54]), .ZN(n3449) );
  NAND2_X1 U3635 ( .A1(n3449), .A2(n3593), .ZN(n3450) );
  NAND2_X1 U3636 ( .A1(p10_C[54]), .A2(n3450), .ZN(n3594) );
  NOR3_X1 U3637 ( .A1(n3590), .A2(n3592), .A3(n3591), .ZN(n3451) );
  NOR2_X1 U3638 ( .A1(p10_S[42]), .A2(p10_C[41]), .ZN(n3452) );
  NAND2_X1 U3639 ( .A1(p10_S[42]), .A2(p10_C[41]), .ZN(n3453) );
  OAI21_X1 U3640 ( .B1(n3451), .B2(n3452), .A(n3453), .ZN(
        p10_Partial_products_sum_add_23_n317) );
  OAI21_X1 U3641 ( .B1(n3573), .B2(n3574), .A(n3575), .ZN(n3454) );
  NAND2_X1 U3642 ( .A1(n3573), .A2(n3574), .ZN(n3455) );
  NAND2_X1 U3643 ( .A1(n3454), .A2(n3455), .ZN(
        p11_Partial_products_sum_add_23_n265) );
  INV_X1 U3644 ( .A(mul4_reg[12]), .ZN(n3456) );
  AOI222_X1 U3645 ( .A1(p9_Partial_products_sum_add_23_n198), .A2(
        p9_Partial_products_sum_add_23_n197), .B1(
        p9_Partial_products_sum_add_23_n198), .B2(
        p9_Partial_products_sum_add_23_n196), .C1(
        p9_Partial_products_sum_add_23_n197), .C2(
        p9_Partial_products_sum_add_23_n196), .ZN(n3457) );
  XOR2_X1 U3646 ( .A(p9_C[54]), .B(p9_final_product2_25_), .Z(n3458) );
  XNOR2_X1 U3647 ( .A(n3457), .B(n3458), .ZN(n3459) );
  INV_X1 U3648 ( .A(n3846), .ZN(n3460) );
  AOI22_X1 U3649 ( .A1(n3846), .A2(n3456), .B1(n3459), .B2(n3460), .ZN(
        REG4_1_n50) );
  INV_X1 U3650 ( .A(reg7[4]), .ZN(n3461) );
  AOI222_X1 U3651 ( .A1(p11_Partial_products_sum_add_23_n285), .A2(
        p11_Partial_products_sum_add_23_n284), .B1(
        p11_Partial_products_sum_add_23_n285), .B2(
        p11_Partial_products_sum_add_23_n283), .C1(
        p11_Partial_products_sum_add_23_n284), .C2(
        p11_Partial_products_sum_add_23_n283), .ZN(n3462) );
  XOR2_X1 U3652 ( .A(p11_S[47]), .B(p11_C[46]), .Z(n3463) );
  XNOR2_X1 U3653 ( .A(n3462), .B(n3463), .ZN(n3464) );
  INV_X1 U3654 ( .A(n3846), .ZN(n3465) );
  AOI22_X1 U3655 ( .A1(n3846), .A2(n3461), .B1(n3464), .B2(n3465), .ZN(
        REG61_n58) );
  OAI21_X1 U3656 ( .B1(p11_Partial_products_sum_add_23_n295), .B2(
        p11_Partial_products_sum_add_23_n296), .A(
        p11_Partial_products_sum_add_23_n297), .ZN(n3559) );
  NAND2_X2 U3657 ( .A1(A1[7]), .A2(n2757), .ZN(n2471) );
  INV_X2 U3658 ( .A(B2[3]), .ZN(n3827) );
  NAND2_X1 U3659 ( .A1(A1[6]), .A2(A1[5]), .ZN(n2472) );
  INV_X2 U3660 ( .A(B2[11]), .ZN(n1085) );
  INV_X2 U3661 ( .A(B2[9]), .ZN(n1104) );
  INV_X1 U3662 ( .A(B2[7]), .ZN(n1118) );
  INV_X2 U3663 ( .A(B2[2]), .ZN(n1234) );
  INV_X2 U3664 ( .A(B3[2]), .ZN(n784) );
  INV_X2 U3665 ( .A(B0[8]), .ZN(n2005) );
  INV_X2 U3666 ( .A(B0[6]), .ZN(n2041) );
  INV_X2 U3667 ( .A(B0[0]), .ZN(n1888) );
  INV_X2 U3668 ( .A(B1[0]), .ZN(n1438) );
  INV_X2 U3669 ( .A(B0[7]), .ZN(n2017) );
  INV_X2 U3670 ( .A(B2[0]), .ZN(n989) );
  INV_X2 U3671 ( .A(B3[0]), .ZN(n539) );
  AND3_X1 U3672 ( .A1(n3601), .A2(n3600), .A3(n3599), .ZN(
        p10_Partial_products_sum_add_23_n283) );
  NAND2_X1 U3673 ( .A1(p6_C[52]), .A2(p6_Partial_products_sum_add_23_n180), 
        .ZN(n3655) );
  AND3_X1 U3674 ( .A1(n3608), .A2(n3607), .A3(n3606), .ZN(
        p10_Partial_products_sum_add_23_n295) );
  AOI222_X2 U3675 ( .A1(p8_S[49]), .A2(p8_C[48]), .B1(p8_S[49]), .B2(n3500), 
        .C1(p8_C[48]), .C2(p8_Partial_products_sum_add_23_n209), .ZN(
        p8_Partial_products_sum_add_23_n205) );
  AOI211_X2 U3676 ( .C1(n3519), .C2(p9_S[45]), .A(n3541), .B(n3534), .ZN(
        p9_Partial_products_sum_add_23_n220) );
  AND2_X1 U3677 ( .A1(p8_Partial_products_sum_add_23_n218), .A2(
        p8_Partial_products_sum_add_23_n219), .ZN(n3512) );
  XNOR2_X1 U3678 ( .A(n1894), .B(n1895), .ZN(p6_S[53]) );
  AOI221_X1 U3679 ( .B1(n2497), .B2(reg2[11]), .C1(n2498), .C2(n3686), .A(
        n2533), .ZN(n2521) );
  AOI221_X1 U3680 ( .B1(n2047), .B2(B0[8]), .C1(n2048), .C2(n2005), .A(n2171), 
        .ZN(n2140) );
  AOI211_X2 U3681 ( .C1(reg1_reg[1]), .C2(reg1_reg[2]), .A(reg1_reg[3]), .B(
        n2322), .ZN(n2148) );
  NAND2_X1 U3682 ( .A1(reg3_reg[1]), .A2(reg3_reg[2]), .ZN(n1213) );
  NAND2_X1 U3683 ( .A1(reg2_reg[1]), .A2(reg2_reg[2]), .ZN(n1662) );
  NAND2_X1 U3684 ( .A1(reg4_reg[1]), .A2(reg4_reg[2]), .ZN(n763) );
  NAND2_X1 U3685 ( .A1(reg1_reg[1]), .A2(reg1_reg[2]), .ZN(n2112) );
  NOR2_X2 U3686 ( .A1(A1[1]), .A2(n2771), .ZN(n2334) );
  INV_X1 U3687 ( .A(B2[6]), .ZN(n1142) );
  NAND2_X1 U3688 ( .A1(A2[7]), .A2(A2[8]), .ZN(n2897) );
  OR2_X1 U3689 ( .A1(A1[6]), .A2(A1[5]), .ZN(n3659) );
  AOI221_X1 U3690 ( .B1(n1878), .B2(B0[0]), .C1(n1879), .C2(n1888), .A(n2207), 
        .ZN(n2194) );
  AOI221_X1 U3691 ( .B1(n1878), .B2(B0[2]), .C1(n1879), .C2(n2133), .A(n2172), 
        .ZN(n2124) );
  AOI221_X1 U3692 ( .B1(n1878), .B2(B0[1]), .C1(n1879), .C2(n1886), .A(n2177), 
        .ZN(n2155) );
  AOI221_X1 U3693 ( .B1(n1878), .B2(B0[6]), .C1(n1879), .C2(n2041), .A(n2062), 
        .ZN(n2061) );
  AOI211_X2 U3694 ( .C1(reg1_reg[11]), .C2(reg1_reg[12]), .A(n2208), .B(n3757), 
        .ZN(n1879) );
  AOI221_X1 U3695 ( .B1(n1428), .B2(B1[0]), .C1(n1429), .C2(n1438), .A(n1757), 
        .ZN(n1744) );
  AOI221_X1 U3696 ( .B1(n1428), .B2(B1[2]), .C1(n1429), .C2(n1683), .A(n1722), 
        .ZN(n1674) );
  AOI221_X1 U3697 ( .B1(n1428), .B2(B1[1]), .C1(n1429), .C2(n1436), .A(n1727), 
        .ZN(n1705) );
  AOI221_X1 U3698 ( .B1(n1428), .B2(B1[6]), .C1(n1429), .C2(n1591), .A(n1612), 
        .ZN(n1611) );
  AOI211_X2 U3699 ( .C1(reg2_reg[11]), .C2(reg2_reg[12]), .A(n1758), .B(n3758), 
        .ZN(n1429) );
  AOI221_X1 U3700 ( .B1(n2328), .B2(reg2[2]), .C1(n2329), .C2(n3692), .A(n2628), .ZN(n2574) );
  AOI221_X1 U3701 ( .B1(n2328), .B2(reg2[0]), .C1(n2329), .C2(n3689), .A(n2660), .ZN(n2647) );
  AOI221_X1 U3702 ( .B1(n2328), .B2(reg2[1]), .C1(n2329), .C2(n3684), .A(n2630), .ZN(n2604) );
  AOI221_X1 U3703 ( .B1(n2328), .B2(reg2[6]), .C1(n2329), .C2(n3687), .A(n2512), .ZN(n2511) );
  AOI211_X2 U3704 ( .C1(A1[11]), .C2(A1[12]), .A(n2661), .B(n2444), .ZN(n2329)
         );
  AOI221_X1 U3705 ( .B1(n979), .B2(B2[0]), .C1(n980), .C2(n989), .A(n1308), 
        .ZN(n1295) );
  AOI221_X1 U3706 ( .B1(n979), .B2(B2[2]), .C1(n980), .C2(n1234), .A(n1273), 
        .ZN(n1225) );
  AOI221_X1 U3707 ( .B1(n979), .B2(B2[1]), .C1(n980), .C2(n987), .A(n1278), 
        .ZN(n1256) );
  AOI221_X1 U3708 ( .B1(n979), .B2(B2[6]), .C1(n980), .C2(n1142), .A(n1163), 
        .ZN(n1162) );
  AOI211_X2 U3709 ( .C1(reg3_reg[11]), .C2(reg3_reg[12]), .A(n1309), .B(n3761), 
        .ZN(n980) );
  AOI221_X1 U3710 ( .B1(n2778), .B2(reg4[0]), .C1(n2779), .C2(n3670), .A(n3106), .ZN(n3093) );
  AOI221_X1 U3711 ( .B1(n2778), .B2(reg4[2]), .C1(n2779), .C2(n3673), .A(n3071), .ZN(n3023) );
  AOI221_X1 U3712 ( .B1(n2778), .B2(reg4[1]), .C1(n2779), .C2(n3666), .A(n3076), .ZN(n3052) );
  AOI221_X1 U3713 ( .B1(n2778), .B2(reg4[6]), .C1(n2779), .C2(n3678), .A(n2962), .ZN(n2961) );
  AOI211_X2 U3714 ( .C1(A2[11]), .C2(A2[12]), .A(n3107), .B(n2894), .ZN(n2779)
         );
  AOI221_X1 U3715 ( .B1(n529), .B2(B3[0]), .C1(n530), .C2(n539), .A(n858), 
        .ZN(n845) );
  AOI221_X1 U3716 ( .B1(n529), .B2(B3[2]), .C1(n530), .C2(n784), .A(n823), 
        .ZN(n775) );
  AOI221_X1 U3717 ( .B1(n529), .B2(B3[1]), .C1(n530), .C2(n537), .A(n828), 
        .ZN(n806) );
  AOI221_X1 U3718 ( .B1(n529), .B2(B3[6]), .C1(n530), .C2(n692), .A(n713), 
        .ZN(n712) );
  AOI211_X2 U3719 ( .C1(reg4_reg[11]), .C2(reg4_reg[12]), .A(n859), .B(n3773), 
        .ZN(n530) );
  AOI221_X1 U3720 ( .B1(n1988), .B2(B0[0]), .C1(n1989), .C2(n1888), .A(n2245), 
        .ZN(n2223) );
  AOI221_X1 U3721 ( .B1(n1988), .B2(B0[2]), .C1(n1989), .C2(n2133), .A(n2222), 
        .ZN(n2196) );
  AOI221_X1 U3722 ( .B1(n1988), .B2(B0[4]), .C1(n1989), .C2(n2075), .A(n2173), 
        .ZN(n2123) );
  AOI221_X1 U3723 ( .B1(n1988), .B2(B0[1]), .C1(n1989), .C2(n1886), .A(n2228), 
        .ZN(n2200) );
  AOI221_X1 U3724 ( .B1(n1988), .B2(B0[5]), .C1(n1989), .C2(n2063), .A(n2143), 
        .ZN(n2117) );
  AOI221_X1 U3725 ( .B1(n1988), .B2(B0[3]), .C1(n1989), .C2(n2115), .A(n2190), 
        .ZN(n2156) );
  AOI211_X4 U3726 ( .C1(reg1_reg[9]), .C2(reg1_reg[10]), .A(reg1_reg[11]), .B(
        n2246), .ZN(n1988) );
  AOI221_X1 U3727 ( .B1(n1538), .B2(B1[0]), .C1(n1539), .C2(n1438), .A(n1795), 
        .ZN(n1773) );
  AOI221_X1 U3728 ( .B1(n1538), .B2(B1[2]), .C1(n1539), .C2(n1683), .A(n1772), 
        .ZN(n1746) );
  AOI221_X1 U3729 ( .B1(n1538), .B2(B1[1]), .C1(n1539), .C2(n1436), .A(n1778), 
        .ZN(n1750) );
  AOI221_X1 U3730 ( .B1(n1538), .B2(B1[4]), .C1(n1539), .C2(n1625), .A(n1723), 
        .ZN(n1673) );
  AOI221_X1 U3731 ( .B1(n1538), .B2(B1[5]), .C1(n1539), .C2(n1613), .A(n1693), 
        .ZN(n1667) );
  AOI221_X1 U3732 ( .B1(n1538), .B2(B1[3]), .C1(n1539), .C2(n1665), .A(n1740), 
        .ZN(n1706) );
  AOI211_X4 U3733 ( .C1(reg2_reg[9]), .C2(reg2_reg[10]), .A(reg2_reg[11]), .B(
        n1796), .ZN(n1538) );
  AOI221_X1 U3734 ( .B1(n1089), .B2(B2[0]), .C1(n1090), .C2(n989), .A(n1345), 
        .ZN(n1323) );
  AOI221_X1 U3735 ( .B1(n1089), .B2(B2[2]), .C1(n1090), .C2(n1234), .A(n1321), 
        .ZN(n1297) );
  AOI221_X1 U3736 ( .B1(n1089), .B2(B2[4]), .C1(n1090), .C2(n1176), .A(n1274), 
        .ZN(n1224) );
  AOI221_X1 U3737 ( .B1(n1089), .B2(B2[1]), .C1(n1090), .C2(n987), .A(n1328), 
        .ZN(n1301) );
  AOI221_X1 U3738 ( .B1(n1089), .B2(B2[5]), .C1(n1090), .C2(n1164), .A(n1244), 
        .ZN(n1218) );
  AOI221_X1 U3739 ( .B1(n1089), .B2(B2[3]), .C1(n1090), .C2(n3827), .A(n1291), 
        .ZN(n1257) );
  AOI211_X4 U3740 ( .C1(reg3_reg[9]), .C2(reg3_reg[10]), .A(reg3_reg[11]), .B(
        n1346), .ZN(n1089) );
  AOI221_X1 U3741 ( .B1(n2888), .B2(reg4[0]), .C1(n2889), .C2(n3670), .A(n3143), .ZN(n3121) );
  AOI221_X1 U3742 ( .B1(n2888), .B2(reg4[4]), .C1(n2889), .C2(n3668), .A(n3072), .ZN(n3022) );
  AOI221_X1 U3743 ( .B1(n2888), .B2(reg4[5]), .C1(n2889), .C2(n3664), .A(n3044), .ZN(n3016) );
  AOI221_X1 U3744 ( .B1(n2888), .B2(reg4[2]), .C1(n2889), .C2(n3673), .A(n3119), .ZN(n3095) );
  AOI221_X1 U3745 ( .B1(n2888), .B2(reg4[1]), .C1(n2889), .C2(n3666), .A(n3126), .ZN(n3099) );
  AOI221_X1 U3746 ( .B1(n2888), .B2(reg4[3]), .C1(n2889), .C2(n3665), .A(n3078), .ZN(n3053) );
  AOI211_X4 U3747 ( .C1(A2[9]), .C2(A2[10]), .A(A2[11]), .B(n3144), .ZN(n2888)
         );
  AOI221_X1 U3748 ( .B1(n639), .B2(B3[0]), .C1(n640), .C2(n539), .A(n896), 
        .ZN(n874) );
  AOI221_X1 U3749 ( .B1(n639), .B2(B3[2]), .C1(n640), .C2(n784), .A(n873), 
        .ZN(n847) );
  AOI221_X1 U3750 ( .B1(n639), .B2(B3[4]), .C1(n640), .C2(n726), .A(n824), 
        .ZN(n774) );
  AOI221_X1 U3751 ( .B1(n639), .B2(B3[5]), .C1(n640), .C2(n714), .A(n794), 
        .ZN(n768) );
  AOI221_X1 U3752 ( .B1(n639), .B2(B3[1]), .C1(n640), .C2(n537), .A(n879), 
        .ZN(n851) );
  AOI221_X1 U3753 ( .B1(n639), .B2(B3[3]), .C1(n640), .C2(n766), .A(n841), 
        .ZN(n807) );
  AOI211_X4 U3754 ( .C1(reg4_reg[9]), .C2(reg4_reg[10]), .A(reg4_reg[11]), .B(
        n897), .ZN(n639) );
  AOI221_X1 U3755 ( .B1(n2006), .B2(B0[4]), .C1(n2007), .C2(n2075), .A(n2212), 
        .ZN(n2192) );
  AOI221_X1 U3756 ( .B1(n2006), .B2(B0[0]), .C1(n2007), .C2(n1888), .A(n2280), 
        .ZN(n2259) );
  AOI221_X1 U3757 ( .B1(n2006), .B2(B0[2]), .C1(n2007), .C2(n2133), .A(n2252), 
        .ZN(n2226) );
  AOI221_X1 U3758 ( .B1(n2006), .B2(B0[3]), .C1(n2007), .C2(n2115), .A(n2230), 
        .ZN(n2199) );
  AOI221_X1 U3759 ( .B1(n2006), .B2(B0[7]), .C1(n2007), .C2(n2017), .A(n2146), 
        .ZN(n2118) );
  AOI221_X1 U3760 ( .B1(n2006), .B2(B0[1]), .C1(n2007), .C2(n1886), .A(n2265), 
        .ZN(n2254) );
  AOI211_X4 U3761 ( .C1(reg1_reg[7]), .C2(reg1_reg[8]), .A(reg1_reg[9]), .B(
        n2281), .ZN(n2006) );
  AOI221_X1 U3762 ( .B1(n1182), .B2(B2[6]), .C1(n1183), .C2(n1142), .A(n1348), 
        .ZN(n1334) );
  AOI221_X1 U3763 ( .B1(n1182), .B2(B2[0]), .C1(n1183), .C2(n989), .A(n1412), 
        .ZN(n1075) );
  AOI221_X1 U3764 ( .B1(n1182), .B2(B2[8]), .C1(n1183), .C2(n1106), .A(n1313), 
        .ZN(n1282) );
  AOI221_X1 U3765 ( .B1(n1182), .B2(B2[5]), .C1(n1183), .C2(n1164), .A(n1372), 
        .ZN(n1357) );
  AOI211_X4 U3766 ( .C1(reg3_reg[3]), .C2(reg3_reg[4]), .A(n3698), .B(n1413), 
        .ZN(n1183) );
  AOI221_X1 U3767 ( .B1(n1631), .B2(B1[0]), .C1(n1632), .C2(n1438), .A(n1862), 
        .ZN(n1524) );
  AOI221_X1 U3768 ( .B1(n1631), .B2(B1[8]), .C1(n1632), .C2(n1555), .A(n1764), 
        .ZN(n1731) );
  AOI221_X1 U3769 ( .B1(n1631), .B2(B1[6]), .C1(n1632), .C2(n1591), .A(n1798), 
        .ZN(n1784) );
  AOI221_X1 U3770 ( .B1(n1631), .B2(B1[7]), .C1(n1632), .C2(n1567), .A(n1790), 
        .ZN(n1771) );
  AOI221_X1 U3771 ( .B1(n1631), .B2(B1[4]), .C1(n1632), .C2(n1625), .A(n1836), 
        .ZN(n1833) );
  AOI211_X4 U3772 ( .C1(reg2_reg[3]), .C2(reg2_reg[4]), .A(n3712), .B(n1863), 
        .ZN(n1632) );
  AOI221_X1 U3773 ( .B1(n732), .B2(B3[0]), .C1(n733), .C2(n539), .A(n963), 
        .ZN(n625) );
  AOI221_X1 U3774 ( .B1(n732), .B2(B3[8]), .C1(n733), .C2(n656), .A(n865), 
        .ZN(n832) );
  AOI221_X1 U3775 ( .B1(n732), .B2(B3[6]), .C1(n733), .C2(n692), .A(n899), 
        .ZN(n885) );
  AOI221_X1 U3776 ( .B1(n732), .B2(B3[4]), .C1(n733), .C2(n726), .A(n937), 
        .ZN(n934) );
  AOI221_X1 U3777 ( .B1(n732), .B2(B3[7]), .C1(n733), .C2(n668), .A(n891), 
        .ZN(n872) );
  AOI211_X4 U3778 ( .C1(reg4_reg[3]), .C2(reg4_reg[4]), .A(n3699), .B(n964), 
        .ZN(n733) );
  AOI221_X1 U3779 ( .B1(n2081), .B2(B0[0]), .C1(n2082), .C2(n1888), .A(n2312), 
        .ZN(n1974) );
  AOI221_X1 U3780 ( .B1(n2081), .B2(B0[6]), .C1(n2082), .C2(n2041), .A(n2248), 
        .ZN(n2234) );
  AOI221_X1 U3781 ( .B1(n2081), .B2(B0[8]), .C1(n2082), .C2(n2005), .A(n2214), 
        .ZN(n2181) );
  AOI221_X1 U3782 ( .B1(n2081), .B2(B0[7]), .C1(n2082), .C2(n2017), .A(n2240), 
        .ZN(n2221) );
  AOI211_X4 U3783 ( .C1(reg1_reg[3]), .C2(reg1_reg[4]), .A(n3711), .B(n2313), 
        .ZN(n2082) );
  AOI221_X1 U3784 ( .B1(n1107), .B2(B2[0]), .C1(n1108), .C2(n989), .A(n1380), 
        .ZN(n1359) );
  AOI221_X1 U3785 ( .B1(n1107), .B2(B2[4]), .C1(n1108), .C2(n1176), .A(n1311), 
        .ZN(n1293) );
  AOI221_X1 U3786 ( .B1(n1107), .B2(B2[2]), .C1(n1108), .C2(n1234), .A(n1352), 
        .ZN(n1326) );
  AOI221_X1 U3787 ( .B1(n1107), .B2(B2[1]), .C1(n1108), .C2(n987), .A(n1365), 
        .ZN(n1354) );
  AOI221_X1 U3788 ( .B1(n1107), .B2(B2[7]), .C1(n1108), .C2(n1118), .A(n1247), 
        .ZN(n1219) );
  AOI211_X4 U3789 ( .C1(reg3_reg[7]), .C2(reg3_reg[8]), .A(reg3_reg[9]), .B(
        n1381), .ZN(n1107) );
  AOI221_X1 U3790 ( .B1(n1556), .B2(B1[0]), .C1(n1557), .C2(n1438), .A(n1830), 
        .ZN(n1809) );
  AOI221_X1 U3791 ( .B1(n1556), .B2(B1[4]), .C1(n1557), .C2(n1625), .A(n1762), 
        .ZN(n1742) );
  AOI221_X1 U3792 ( .B1(n1556), .B2(B1[2]), .C1(n1557), .C2(n1683), .A(n1802), 
        .ZN(n1776) );
  AOI221_X1 U3793 ( .B1(n1556), .B2(B1[7]), .C1(n1557), .C2(n1567), .A(n1696), 
        .ZN(n1668) );
  AOI221_X1 U3794 ( .B1(n1556), .B2(B1[1]), .C1(n1557), .C2(n1436), .A(n1815), 
        .ZN(n1804) );
  AOI211_X4 U3795 ( .C1(reg2_reg[7]), .C2(reg2_reg[8]), .A(reg2_reg[9]), .B(
        n1831), .ZN(n1556) );
  AOI221_X1 U3796 ( .B1(n657), .B2(B3[0]), .C1(n658), .C2(n539), .A(n931), 
        .ZN(n910) );
  AOI221_X1 U3797 ( .B1(n657), .B2(B3[4]), .C1(n658), .C2(n726), .A(n863), 
        .ZN(n843) );
  AOI221_X1 U3798 ( .B1(n657), .B2(B3[2]), .C1(n658), .C2(n784), .A(n903), 
        .ZN(n877) );
  AOI221_X1 U3799 ( .B1(n657), .B2(B3[1]), .C1(n658), .C2(n537), .A(n916), 
        .ZN(n905) );
  AOI221_X1 U3800 ( .B1(n657), .B2(B3[7]), .C1(n658), .C2(n668), .A(n797), 
        .ZN(n769) );
  AOI211_X4 U3801 ( .C1(reg4_reg[7]), .C2(reg4_reg[8]), .A(reg4_reg[9]), .B(
        n932), .ZN(n657) );
  AOI211_X4 U3802 ( .C1(A1[9]), .C2(A1[10]), .A(A1[11]), .B(n2698), .ZN(n2438)
         );
  AOI211_X4 U3803 ( .C1(reg1_reg[6]), .C2(reg1_reg[5]), .A(reg1_reg[7]), .B(
        n2304), .ZN(n2047) );
  AOI221_X1 U3804 ( .B1(n1597), .B2(B1[4]), .C1(n1598), .C2(n1625), .A(n1799), 
        .ZN(n1783) );
  AOI221_X1 U3805 ( .B1(n1597), .B2(B1[2]), .C1(n1598), .C2(n1683), .A(n1832), 
        .ZN(n1812) );
  AOI221_X1 U3806 ( .B1(n1597), .B2(B1[3]), .C1(n1598), .C2(n1665), .A(n1823), 
        .ZN(n1803) );
  AOI221_X1 U3807 ( .B1(n1597), .B2(B1[8]), .C1(n1598), .C2(n1555), .A(n1721), 
        .ZN(n1690) );
  AOI211_X4 U3808 ( .C1(reg2_reg[5]), .C2(reg2_reg[6]), .A(n3714), .B(n1854), 
        .ZN(n1598) );
  AOI221_X1 U3809 ( .B1(n698), .B2(B3[4]), .C1(n699), .C2(n726), .A(n900), 
        .ZN(n884) );
  AOI221_X1 U3810 ( .B1(n698), .B2(B3[2]), .C1(n699), .C2(n784), .A(n933), 
        .ZN(n913) );
  AOI221_X1 U3811 ( .B1(n698), .B2(B3[3]), .C1(n699), .C2(n766), .A(n924), 
        .ZN(n904) );
  AOI221_X1 U3812 ( .B1(n698), .B2(B3[8]), .C1(n699), .C2(n656), .A(n822), 
        .ZN(n791) );
  AOI211_X4 U3813 ( .C1(reg4_reg[5]), .C2(reg4_reg[6]), .A(n3697), .B(n955), 
        .ZN(n699) );
  AOI211_X4 U3814 ( .C1(reg1_reg[7]), .C2(reg1_reg[8]), .A(n3713), .B(n2281), 
        .ZN(n2007) );
  AOI211_X4 U3815 ( .C1(reg3_reg[7]), .C2(reg3_reg[8]), .A(n3721), .B(n1381), 
        .ZN(n1108) );
  AOI211_X4 U3816 ( .C1(reg2_reg[7]), .C2(reg2_reg[8]), .A(n3719), .B(n1831), 
        .ZN(n1557) );
  AOI211_X4 U3817 ( .C1(reg4_reg[7]), .C2(reg4_reg[8]), .A(n3720), .B(n932), 
        .ZN(n658) );
  AOI211_X4 U3818 ( .C1(reg1_reg[9]), .C2(reg1_reg[10]), .A(n3674), .B(n2246), 
        .ZN(n1989) );
  AOI211_X4 U3819 ( .C1(reg3_reg[9]), .C2(reg3_reg[10]), .A(n3695), .B(n1346), 
        .ZN(n1090) );
  AOI211_X4 U3820 ( .C1(reg2_reg[9]), .C2(reg2_reg[10]), .A(n3694), .B(n1796), 
        .ZN(n1539) );
  AOI211_X4 U3821 ( .C1(reg4_reg[9]), .C2(reg4_reg[10]), .A(n3675), .B(n897), 
        .ZN(n640) );
  AOI211_X4 U3822 ( .C1(A2[9]), .C2(A2[10]), .A(n3120), .B(n3144), .ZN(n2889)
         );
  AOI211_X4 U3823 ( .C1(reg1_reg[5]), .C2(reg1_reg[6]), .A(n3710), .B(n2304), 
        .ZN(n2048) );
  AOI211_X4 U3824 ( .C1(A2[12]), .C2(A2[11]), .A(A2[13]), .B(n3107), .ZN(n2778) );
  AOI211_X4 U3825 ( .C1(A1[12]), .C2(A1[11]), .A(A1[13]), .B(n2661), .ZN(n2328) );
  AOI211_X4 U3826 ( .C1(reg3_reg[3]), .C2(reg3_reg[4]), .A(reg3_reg[5]), .B(
        n1413), .ZN(n1182) );
  AOI211_X4 U3827 ( .C1(reg4_reg[3]), .C2(reg4_reg[4]), .A(reg4_reg[5]), .B(
        n964), .ZN(n732) );
  AOI211_X4 U3828 ( .C1(reg2_reg[3]), .C2(reg2_reg[4]), .A(reg2_reg[5]), .B(
        n1863), .ZN(n1631) );
  AOI222_X4 U3829 ( .A1(n1931), .A2(n1932), .B1(n1931), .B2(n1929), .C1(n1932), 
        .C2(n1929), .ZN(p6_C[44]) );
  NOR2_X2 U3830 ( .A1(A2[1]), .A2(n3218), .ZN(n2784) );
  AOI211_X4 U3831 ( .C1(reg3_reg[6]), .C2(reg3_reg[5]), .A(reg3_reg[7]), .B(
        n1404), .ZN(n1148) );
  AOI211_X4 U3832 ( .C1(reg4_reg[6]), .C2(reg4_reg[5]), .A(reg4_reg[7]), .B(
        n955), .ZN(n698) );
  AOI211_X4 U3833 ( .C1(reg2_reg[6]), .C2(reg2_reg[5]), .A(reg2_reg[7]), .B(
        n1854), .ZN(n1597) );
  AOI211_X4 U3834 ( .C1(reg3_reg[1]), .C2(reg3_reg[2]), .A(n3702), .B(n1422), 
        .ZN(n1250) );
  AOI211_X4 U3835 ( .C1(A1[9]), .C2(A1[10]), .A(n2674), .B(n2698), .ZN(n2439)
         );
  AOI211_X4 U3836 ( .C1(reg4_reg[12]), .C2(reg4_reg[11]), .A(reg4_reg[13]), 
        .B(n859), .ZN(n529) );
  AOI211_X4 U3837 ( .C1(reg2_reg[12]), .C2(reg2_reg[11]), .A(reg2_reg[13]), 
        .B(n1758), .ZN(n1428) );
  AOI211_X4 U3838 ( .C1(reg3_reg[12]), .C2(reg3_reg[11]), .A(reg3_reg[13]), 
        .B(n1309), .ZN(n979) );
  AOI211_X4 U3839 ( .C1(reg1_reg[12]), .C2(reg1_reg[11]), .A(reg1_reg[13]), 
        .B(n2208), .ZN(n1878) );
  AOI211_X4 U3840 ( .C1(reg1_reg[3]), .C2(reg1_reg[4]), .A(reg1_reg[5]), .B(
        n2313), .ZN(n2081) );
  AOI211_X4 U3841 ( .C1(reg4_reg[1]), .C2(reg4_reg[2]), .A(reg4_reg[3]), .B(
        n973), .ZN(n799) );
  AOI211_X4 U3842 ( .C1(reg2_reg[1]), .C2(reg2_reg[2]), .A(reg2_reg[3]), .B(
        n1872), .ZN(n1698) );
  OAI21_X1 U3843 ( .B1(p7_Partial_products_sum_add_23_n241), .B2(
        p7_Partial_products_sum_add_23_n242), .A(
        p7_Partial_products_sum_add_23_n243), .ZN(
        p7_Partial_products_sum_add_23_n240) );
  XNOR2_X1 U3844 ( .A(n3481), .B(p7_Partial_products_sum_add_23_n216), .ZN(
        temp2[4]) );
  XNOR2_X1 U3845 ( .A(p7_Partial_products_sum_add_23_n198), .B(n3495), .ZN(
        temp2[10]) );
  XNOR2_X1 U3846 ( .A(p7_Partial_products_sum_add_23_n204), .B(
        p7_Partial_products_sum_add_23_n203), .ZN(temp2[8]) );
  XNOR2_X1 U3847 ( .A(p7_Partial_products_sum_add_23_n222), .B(n3493), .ZN(
        temp2[2]) );
  OAI21_X1 U3848 ( .B1(p7_Partial_products_sum_add_23_n237), .B2(
        p7_Partial_products_sum_add_23_n238), .A(
        p7_Partial_products_sum_add_23_n239), .ZN(
        p7_Partial_products_sum_add_23_n236) );
  XNOR2_X1 U3849 ( .A(n3497), .B(p7_Partial_products_sum_add_23_n192), .ZN(
        temp2[12]) );
  XNOR2_X1 U3850 ( .A(p7_Partial_products_sum_add_23_n210), .B(n3488), .ZN(
        temp2[6]) );
  XNOR2_X1 U3851 ( .A(p7_Partial_products_sum_add_23_n189), .B(
        p7_Partial_products_sum_add_23_n190), .ZN(temp2[13]) );
  OAI21_X1 U3852 ( .B1(p7_Partial_products_sum_add_23_n229), .B2(
        p7_Partial_products_sum_add_23_n230), .A(
        p7_Partial_products_sum_add_23_n231), .ZN(
        p7_Partial_products_sum_add_23_n227) );
  NAND2_X1 U3853 ( .A1(p7_Partial_products_sum_add_23_n249), .A2(
        p7_Partial_products_sum_add_23_n250), .ZN(
        p7_Partial_products_sum_add_23_n248) );
  AOI222_X1 U3854 ( .A1(p7_Partial_products_sum_add_23_n217), .A2(
        p7_Partial_products_sum_add_23_n218), .B1(
        p7_Partial_products_sum_add_23_n217), .B2(
        p7_Partial_products_sum_add_23_n219), .C1(
        p7_Partial_products_sum_add_23_n218), .C2(
        p7_Partial_products_sum_add_23_n219), .ZN(
        p7_Partial_products_sum_add_23_n215) );
  AOI222_X1 U3855 ( .A1(p7_Partial_products_sum_add_23_n211), .A2(
        p7_Partial_products_sum_add_23_n212), .B1(
        p7_Partial_products_sum_add_23_n211), .B2(
        p7_Partial_products_sum_add_23_n213), .C1(
        p7_Partial_products_sum_add_23_n212), .C2(
        p7_Partial_products_sum_add_23_n213), .ZN(
        p7_Partial_products_sum_add_23_n209) );
  AOI222_X1 U3856 ( .A1(p7_Partial_products_sum_add_23_n211), .A2(
        p7_Partial_products_sum_add_23_n212), .B1(
        p7_Partial_products_sum_add_23_n211), .B2(
        p7_Partial_products_sum_add_23_n213), .C1(
        p7_Partial_products_sum_add_23_n212), .C2(
        p7_Partial_products_sum_add_23_n213), .ZN(n3482) );
  NOR3_X1 U3857 ( .A1(n3485), .A2(n3484), .A3(n3483), .ZN(
        p7_Partial_products_sum_add_23_n189) );
  NAND2_X1 U3858 ( .A1(p7_S[35]), .A2(p7_C[34]), .ZN(n3486) );
  NAND2_X1 U3859 ( .A1(p7_Partial_products_sum_add_23_n240), .A2(p7_C[36]), 
        .ZN(n3487) );
  OAI21_X1 U3860 ( .B1(p7_Partial_products_sum_add_23_n233), .B2(
        p7_Partial_products_sum_add_23_n234), .A(
        p7_Partial_products_sum_add_23_n235), .ZN(
        p7_Partial_products_sum_add_23_n232) );
  XNOR2_X1 U3861 ( .A(p7_Partial_products_sum_add_23_n205), .B(
        p7_Partial_products_sum_add_23_n208), .ZN(temp2[7]) );
  NAND2_X1 U3862 ( .A1(p7_Partial_products_sum_add_23_n236), .A2(p7_C[38]), 
        .ZN(n3489) );
  NAND2_X1 U3863 ( .A1(p7_C[48]), .A2(p7_Partial_products_sum_add_23_n209), 
        .ZN(n3490) );
  NAND2_X1 U3864 ( .A1(p7_S[49]), .A2(n3482), .ZN(n3491) );
  NAND2_X1 U3865 ( .A1(p7_S[49]), .A2(p7_C[48]), .ZN(n3492) );
  NOR2_X1 U3866 ( .A1(p7_C[41]), .A2(p7_S[42]), .ZN(
        p7_Partial_products_sum_add_23_n230) );
  NAND2_X1 U3867 ( .A1(p7_C[41]), .A2(p7_S[42]), .ZN(
        p7_Partial_products_sum_add_23_n231) );
  AOI222_X1 U3868 ( .A1(p7_Partial_products_sum_add_23_n223), .A2(
        p7_Partial_products_sum_add_23_n224), .B1(
        p7_Partial_products_sum_add_23_n223), .B2(
        p7_Partial_products_sum_add_23_n225), .C1(
        p7_Partial_products_sum_add_23_n224), .C2(
        p7_Partial_products_sum_add_23_n225), .ZN(
        p7_Partial_products_sum_add_23_n221) );
  AOI222_X1 U3869 ( .A1(p7_Partial_products_sum_add_23_n199), .A2(
        p7_Partial_products_sum_add_23_n200), .B1(
        p7_Partial_products_sum_add_23_n199), .B2(
        p7_Partial_products_sum_add_23_n201), .C1(
        p7_Partial_products_sum_add_23_n200), .C2(
        p7_Partial_products_sum_add_23_n201), .ZN(
        p7_Partial_products_sum_add_23_n197) );
  AOI222_X1 U3870 ( .A1(p7_Partial_products_sum_add_23_n193), .A2(
        p7_Partial_products_sum_add_23_n194), .B1(
        p7_Partial_products_sum_add_23_n193), .B2(
        p7_Partial_products_sum_add_23_n195), .C1(
        p7_Partial_products_sum_add_23_n194), .C2(
        p7_Partial_products_sum_add_23_n195), .ZN(
        p7_Partial_products_sum_add_23_n191) );
  AOI222_X1 U3871 ( .A1(p7_Partial_products_sum_add_23_n223), .A2(
        p7_Partial_products_sum_add_23_n224), .B1(
        p7_Partial_products_sum_add_23_n223), .B2(
        p7_Partial_products_sum_add_23_n225), .C1(
        p7_Partial_products_sum_add_23_n224), .C2(
        p7_Partial_products_sum_add_23_n225), .ZN(n3494) );
  AOI222_X1 U3872 ( .A1(p7_Partial_products_sum_add_23_n199), .A2(
        p7_Partial_products_sum_add_23_n200), .B1(
        p7_Partial_products_sum_add_23_n199), .B2(
        p7_Partial_products_sum_add_23_n201), .C1(
        p7_Partial_products_sum_add_23_n200), .C2(
        p7_Partial_products_sum_add_23_n201), .ZN(n3496) );
  AOI222_X1 U3873 ( .A1(p7_Partial_products_sum_add_23_n193), .A2(
        p7_Partial_products_sum_add_23_n194), .B1(
        p7_Partial_products_sum_add_23_n193), .B2(
        p7_Partial_products_sum_add_23_n195), .C1(
        p7_Partial_products_sum_add_23_n194), .C2(
        p7_Partial_products_sum_add_23_n195), .ZN(n3498) );
  AOI222_X1 U3874 ( .A1(p7_Partial_products_sum_add_23_n232), .A2(p7_S[41]), 
        .B1(p7_Partial_products_sum_add_23_n232), .B2(p7_C[40]), .C1(p7_S[41]), 
        .C2(p7_C[40]), .ZN(p7_Partial_products_sum_add_23_n229) );
  AOI222_X1 U3875 ( .A1(p7_Partial_products_sum_add_23_n193), .A2(
        p7_Partial_products_sum_add_23_n194), .B1(
        p7_Partial_products_sum_add_23_n193), .B2(
        p7_Partial_products_sum_add_23_n195), .C1(
        p7_Partial_products_sum_add_23_n194), .C2(
        p7_Partial_products_sum_add_23_n195), .ZN(n3497) );
  AOI222_X1 U3876 ( .A1(p7_Partial_products_sum_add_23_n217), .A2(
        p7_Partial_products_sum_add_23_n218), .B1(
        p7_Partial_products_sum_add_23_n217), .B2(
        p7_Partial_products_sum_add_23_n219), .C1(
        p7_Partial_products_sum_add_23_n218), .C2(
        p7_Partial_products_sum_add_23_n219), .ZN(n3481) );
  AOI222_X1 U3877 ( .A1(p7_Partial_products_sum_add_23_n199), .A2(
        p7_Partial_products_sum_add_23_n200), .B1(
        p7_Partial_products_sum_add_23_n199), .B2(
        p7_Partial_products_sum_add_23_n201), .C1(
        p7_Partial_products_sum_add_23_n200), .C2(
        p7_Partial_products_sum_add_23_n201), .ZN(n3495) );
  AOI222_X1 U3878 ( .A1(p7_Partial_products_sum_add_23_n211), .A2(
        p7_Partial_products_sum_add_23_n212), .B1(
        p7_Partial_products_sum_add_23_n211), .B2(
        p7_Partial_products_sum_add_23_n213), .C1(
        p7_Partial_products_sum_add_23_n212), .C2(
        p7_Partial_products_sum_add_23_n213), .ZN(n3488) );
  AOI222_X1 U3879 ( .A1(p7_Partial_products_sum_add_23_n223), .A2(
        p7_Partial_products_sum_add_23_n224), .B1(
        p7_Partial_products_sum_add_23_n223), .B2(
        p7_Partial_products_sum_add_23_n225), .C1(
        p7_Partial_products_sum_add_23_n224), .C2(
        p7_Partial_products_sum_add_23_n225), .ZN(n3493) );
  AND2_X1 U3880 ( .A1(p7_C[54]), .A2(p7_final_product2_25_), .ZN(n3485) );
  AND3_X1 U3881 ( .A1(p7_final_product1[0]), .A2(reg2_reg[1]), .A3(
        p7_final_product1[1]), .ZN(n3499) );
  AOI222_X1 U3882 ( .A1(p7_Partial_products_sum_add_23_n205), .A2(
        p7_Partial_products_sum_add_23_n206), .B1(
        p7_Partial_products_sum_add_23_n205), .B2(
        p7_Partial_products_sum_add_23_n207), .C1(
        p7_Partial_products_sum_add_23_n206), .C2(
        p7_Partial_products_sum_add_23_n207), .ZN(
        p7_Partial_products_sum_add_23_n203) );
  AND2_X1 U3883 ( .A1(p7_C[54]), .A2(n3498), .ZN(n3484) );
  AND2_X1 U3884 ( .A1(p7_final_product2_25_), .A2(
        p7_Partial_products_sum_add_23_n191), .ZN(n3483) );
  AOI222_X4 U3885 ( .A1(p7_S[43]), .A2(p7_C[42]), .B1(p7_S[43]), .B2(
        p7_Partial_products_sum_add_23_n227), .C1(p7_C[42]), .C2(
        p7_Partial_products_sum_add_23_n227), .ZN(
        p7_Partial_products_sum_add_23_n223) );
  AOI222_X4 U3886 ( .A1(p7_S[51]), .A2(p7_C[50]), .B1(p7_S[51]), .B2(
        p7_Partial_products_sum_add_23_n203), .C1(p7_C[50]), .C2(
        p7_Partial_products_sum_add_23_n203), .ZN(
        p7_Partial_products_sum_add_23_n199) );
  AOI222_X4 U3887 ( .A1(p7_S[47]), .A2(p7_C[46]), .B1(p7_S[47]), .B2(n3481), 
        .C1(p7_C[46]), .C2(p7_Partial_products_sum_add_23_n215), .ZN(
        p7_Partial_products_sum_add_23_n211) );
  AOI222_X4 U3888 ( .A1(p7_S[53]), .A2(p7_C[52]), .B1(p7_S[53]), .B2(n3496), 
        .C1(p7_C[52]), .C2(p7_Partial_products_sum_add_23_n197), .ZN(
        p7_Partial_products_sum_add_23_n193) );
  AND3_X2 U3889 ( .A1(n3492), .A2(n3491), .A3(n3490), .ZN(
        p7_Partial_products_sum_add_23_n205) );
  AOI222_X4 U3890 ( .A1(p7_S[45]), .A2(p7_C[44]), .B1(p7_S[45]), .B2(n3494), 
        .C1(p7_C[44]), .C2(p7_Partial_products_sum_add_23_n221), .ZN(
        p7_Partial_products_sum_add_23_n217) );
  AOI222_X1 U3891 ( .A1(p8_Partial_products_sum_add_23_n211), .A2(
        p8_Partial_products_sum_add_23_n212), .B1(
        p8_Partial_products_sum_add_23_n211), .B2(
        p8_Partial_products_sum_add_23_n213), .C1(
        p8_Partial_products_sum_add_23_n212), .C2(
        p8_Partial_products_sum_add_23_n213), .ZN(
        p8_Partial_products_sum_add_23_n209) );
  OAI21_X1 U3892 ( .B1(p8_Partial_products_sum_add_23_n245), .B2(
        p8_Partial_products_sum_add_23_n246), .A(
        p8_Partial_products_sum_add_23_n247), .ZN(
        p8_Partial_products_sum_add_23_n244) );
  OAI21_X1 U3893 ( .B1(p8_Partial_products_sum_add_23_n241), .B2(
        p8_Partial_products_sum_add_23_n242), .A(
        p8_Partial_products_sum_add_23_n243), .ZN(
        p8_Partial_products_sum_add_23_n240) );
  XNOR2_X1 U3894 ( .A(p8_Partial_products_sum_add_23_n210), .B(n3500), .ZN(
        temp3[6]) );
  XNOR2_X1 U3895 ( .A(p8_Partial_products_sum_add_23_n204), .B(
        p8_Partial_products_sum_add_23_n203), .ZN(temp3[8]) );
  XNOR2_X1 U3896 ( .A(p8_Partial_products_sum_add_23_n222), .B(
        p8_Partial_products_sum_add_23_n221), .ZN(temp3[2]) );
  OAI21_X1 U3897 ( .B1(p8_Partial_products_sum_add_23_n237), .B2(
        p8_Partial_products_sum_add_23_n238), .A(
        p8_Partial_products_sum_add_23_n239), .ZN(
        p8_Partial_products_sum_add_23_n236) );
  NAND2_X1 U3898 ( .A1(p8_S[35]), .A2(p8_C[34]), .ZN(n3501) );
  NAND2_X1 U3899 ( .A1(p8_Partial_products_sum_add_23_n240), .A2(p8_C[36]), 
        .ZN(n3502) );
  NOR2_X1 U3900 ( .A1(p8_S[42]), .A2(p8_C[41]), .ZN(
        p8_Partial_products_sum_add_23_n230) );
  NAND2_X1 U3901 ( .A1(p8_C[41]), .A2(p8_S[42]), .ZN(
        p8_Partial_products_sum_add_23_n231) );
  XNOR2_X1 U3902 ( .A(p8_Partial_products_sum_add_23_n198), .B(
        p8_Partial_products_sum_add_23_n197), .ZN(temp3[10]) );
  XNOR2_X1 U3903 ( .A(p8_Partial_products_sum_add_23_n205), .B(
        p8_Partial_products_sum_add_23_n208), .ZN(temp3[7]) );
  OAI21_X1 U3904 ( .B1(p8_Partial_products_sum_add_23_n233), .B2(
        p8_Partial_products_sum_add_23_n234), .A(
        p8_Partial_products_sum_add_23_n235), .ZN(
        p8_Partial_products_sum_add_23_n232) );
  XNOR2_X1 U3905 ( .A(p8_Partial_products_sum_add_23_n216), .B(
        p8_Partial_products_sum_add_23_n215), .ZN(temp3[4]) );
  AOI222_X1 U3906 ( .A1(p8_Partial_products_sum_add_23_n236), .A2(p8_S[39]), 
        .B1(p8_Partial_products_sum_add_23_n236), .B2(p8_C[38]), .C1(p8_S[39]), 
        .C2(p8_C[38]), .ZN(p8_Partial_products_sum_add_23_n233) );
  NAND2_X1 U3907 ( .A1(p8_Partial_products_sum_add_23_n249), .A2(
        p8_Partial_products_sum_add_23_n250), .ZN(
        p8_Partial_products_sum_add_23_n248) );
  AOI222_X1 U3908 ( .A1(p8_S[33]), .A2(p8_C[32]), .B1(p8_S[33]), .B2(
        p8_Partial_products_sum_add_23_n248), .C1(p8_C[32]), .C2(
        p8_Partial_products_sum_add_23_n248), .ZN(
        p8_Partial_products_sum_add_23_n245) );
  OAI21_X1 U3909 ( .B1(p8_Partial_products_sum_add_23_n229), .B2(
        p8_Partial_products_sum_add_23_n230), .A(
        p8_Partial_products_sum_add_23_n231), .ZN(
        p8_Partial_products_sum_add_23_n227) );
  XNOR2_X1 U3910 ( .A(p8_Partial_products_sum_add_23_n228), .B(
        p8_Partial_products_sum_add_23_n227), .ZN(temp3[0]) );
  XNOR2_X1 U3911 ( .A(p8_Partial_products_sum_add_23_n223), .B(
        p8_Partial_products_sum_add_23_n226), .ZN(temp3[1]) );
  NOR2_X1 U3912 ( .A1(p8_S[34]), .A2(p8_C[33]), .ZN(
        p8_Partial_products_sum_add_23_n246) );
  XNOR2_X1 U3913 ( .A(p8_Partial_products_sum_add_23_n193), .B(
        p8_Partial_products_sum_add_23_n196), .ZN(temp3[11]) );
  AOI222_X1 U3914 ( .A1(p8_Partial_products_sum_add_23_n211), .A2(
        p8_Partial_products_sum_add_23_n212), .B1(
        p8_Partial_products_sum_add_23_n211), .B2(
        p8_Partial_products_sum_add_23_n213), .C1(
        p8_Partial_products_sum_add_23_n212), .C2(
        p8_Partial_products_sum_add_23_n213), .ZN(n3500) );
  AOI22_X1 U3915 ( .A1(p8_S[44]), .A2(p8_C[43]), .B1(
        p8_Partial_products_sum_add_23_n225), .B2(
        p8_Partial_products_sum_add_23_n224), .ZN(
        p8_Partial_products_sum_add_23_n226) );
  NAND2_X1 U3916 ( .A1(p8_Partial_products_sum_add_23_n232), .A2(p8_C[40]), 
        .ZN(n3503) );
  XNOR2_X1 U3917 ( .A(p8_Partial_products_sum_add_23_n189), .B(
        p8_Partial_products_sum_add_23_n190), .ZN(temp3[13]) );
  NAND2_X1 U3918 ( .A1(p8_C[54]), .A2(p8_Partial_products_sum_add_23_n191), 
        .ZN(n3505) );
  AOI222_X1 U3919 ( .A1(p8_Partial_products_sum_add_23_n193), .A2(
        p8_Partial_products_sum_add_23_n194), .B1(
        p8_Partial_products_sum_add_23_n193), .B2(
        p8_Partial_products_sum_add_23_n195), .C1(
        p8_Partial_products_sum_add_23_n194), .C2(
        p8_Partial_products_sum_add_23_n195), .ZN(n3504) );
  AOI222_X1 U3920 ( .A1(p8_Partial_products_sum_add_23_n193), .A2(
        p8_Partial_products_sum_add_23_n194), .B1(
        p8_Partial_products_sum_add_23_n193), .B2(
        p8_Partial_products_sum_add_23_n195), .C1(
        p8_Partial_products_sum_add_23_n194), .C2(
        p8_Partial_products_sum_add_23_n195), .ZN(
        p8_Partial_products_sum_add_23_n191) );
  NAND2_X1 U3921 ( .A1(p8_Partial_products_sum_add_23_n197), .A2(p8_S[53]), 
        .ZN(n3507) );
  NAND2_X1 U3922 ( .A1(p8_Partial_products_sum_add_23_n197), .A2(p8_C[52]), 
        .ZN(n3508) );
  OAI21_X1 U3923 ( .B1(p8_Partial_products_sum_add_23_n201), .B2(
        p8_Partial_products_sum_add_23_n200), .A(
        p8_Partial_products_sum_add_23_n199), .ZN(n3510) );
  AOI222_X1 U3924 ( .A1(p8_S[45]), .A2(p8_C[44]), .B1(p8_S[45]), .B2(
        p8_Partial_products_sum_add_23_n221), .C1(p8_C[44]), .C2(
        p8_Partial_products_sum_add_23_n221), .ZN(
        p8_Partial_products_sum_add_23_n217) );
  NAND2_X1 U3925 ( .A1(p8_Partial_products_sum_add_23_n201), .A2(
        p8_Partial_products_sum_add_23_n200), .ZN(n3509) );
  NAND2_X1 U3926 ( .A1(p8_S[53]), .A2(p8_C[52]), .ZN(n3506) );
  INV_X1 U3927 ( .A(p8_S[44]), .ZN(p8_Partial_products_sum_add_23_n224) );
  AND2_X1 U3928 ( .A1(n3510), .A2(n3509), .ZN(
        p8_Partial_products_sum_add_23_n197) );
  AOI222_X4 U3929 ( .A1(p8_S[47]), .A2(p8_C[46]), .B1(p8_S[47]), .B2(
        p8_Partial_products_sum_add_23_n215), .C1(p8_C[46]), .C2(
        p8_Partial_products_sum_add_23_n215), .ZN(
        p8_Partial_products_sum_add_23_n211) );
  AOI222_X4 U3930 ( .A1(p8_S[43]), .A2(p8_C[42]), .B1(p8_S[43]), .B2(
        p8_Partial_products_sum_add_23_n227), .C1(p8_C[42]), .C2(
        p8_Partial_products_sum_add_23_n227), .ZN(
        p8_Partial_products_sum_add_23_n223) );
  AND3_X2 U3931 ( .A1(n3508), .A2(n3507), .A3(n3506), .ZN(
        p8_Partial_products_sum_add_23_n193) );
  NOR3_X1 U3932 ( .A1(n3514), .A2(n3513), .A3(n3512), .ZN(
        p8_Partial_products_sum_add_23_n215) );
  AND2_X1 U3933 ( .A1(p8_Partial_products_sum_add_23_n217), .A2(
        p8_Partial_products_sum_add_23_n219), .ZN(n3513) );
  AND2_X1 U3934 ( .A1(p8_Partial_products_sum_add_23_n217), .A2(
        p8_Partial_products_sum_add_23_n218), .ZN(n3514) );
  NAND2_X1 U3935 ( .A1(p8_Partial_products_sum_add_23_n205), .A2(
        p8_Partial_products_sum_add_23_n207), .ZN(n3515) );
  NOR3_X1 U3936 ( .A1(n3518), .A2(n3517), .A3(n3516), .ZN(
        p8_Partial_products_sum_add_23_n199) );
  AND2_X1 U3937 ( .A1(p8_C[50]), .A2(p8_Partial_products_sum_add_23_n203), 
        .ZN(n3516) );
  AND2_X1 U3938 ( .A1(p8_S[51]), .A2(p8_Partial_products_sum_add_23_n203), 
        .ZN(n3517) );
  AND2_X1 U3939 ( .A1(p8_S[51]), .A2(p8_C[50]), .ZN(n3518) );
  OAI21_X1 U3940 ( .B1(p9_Partial_products_sum_add_23_n244), .B2(
        p9_Partial_products_sum_add_23_n245), .A(
        p9_Partial_products_sum_add_23_n246), .ZN(
        p9_Partial_products_sum_add_23_n243) );
  XNOR2_X1 U3941 ( .A(p9_Partial_products_sum_add_23_n219), .B(n3521), .ZN(
        temp4[4]) );
  XNOR2_X1 U3942 ( .A(p9_Partial_products_sum_add_23_n201), .B(n3522), .ZN(
        temp4[10]) );
  XNOR2_X1 U3943 ( .A(p9_Partial_products_sum_add_23_n207), .B(n3520), .ZN(
        temp4[8]) );
  XNOR2_X1 U3944 ( .A(p9_Partial_products_sum_add_23_n225), .B(n3519), .ZN(
        temp4[2]) );
  OAI21_X1 U3945 ( .B1(p9_Partial_products_sum_add_23_n248), .B2(
        p9_Partial_products_sum_add_23_n249), .A(
        p9_Partial_products_sum_add_23_n250), .ZN(
        p9_Partial_products_sum_add_23_n247) );
  OAI21_X1 U3946 ( .B1(p9_Partial_products_sum_add_23_n240), .B2(
        p9_Partial_products_sum_add_23_n241), .A(
        p9_Partial_products_sum_add_23_n242), .ZN(
        p9_Partial_products_sum_add_23_n239) );
  XNOR2_X1 U3947 ( .A(p9_Partial_products_sum_add_23_n208), .B(
        p9_Partial_products_sum_add_23_n211), .ZN(temp4[7]) );
  XNOR2_X1 U3948 ( .A(p9_Partial_products_sum_add_23_n226), .B(
        p9_Partial_products_sum_add_23_n229), .ZN(temp4[1]) );
  XNOR2_X1 U3949 ( .A(p9_Partial_products_sum_add_23_n213), .B(n3525), .ZN(
        temp4[6]) );
  AOI222_X1 U3950 ( .A1(p9_Partial_products_sum_add_23_n220), .A2(
        p9_Partial_products_sum_add_23_n221), .B1(
        p9_Partial_products_sum_add_23_n220), .B2(
        p9_Partial_products_sum_add_23_n222), .C1(
        p9_Partial_products_sum_add_23_n221), .C2(
        p9_Partial_products_sum_add_23_n222), .ZN(n3521) );
  NAND2_X1 U3951 ( .A1(p9_S[35]), .A2(p9_C[34]), .ZN(n3523) );
  NAND2_X1 U3952 ( .A1(p9_Partial_products_sum_add_23_n243), .A2(p9_C[36]), 
        .ZN(n3524) );
  AOI222_X1 U3953 ( .A1(p9_Partial_products_sum_add_23_n239), .A2(p9_S[39]), 
        .B1(p9_Partial_products_sum_add_23_n239), .B2(p9_C[38]), .C1(p9_S[39]), 
        .C2(p9_C[38]), .ZN(p9_Partial_products_sum_add_23_n236) );
  AOI222_X1 U3954 ( .A1(p9_S[33]), .A2(p9_C[32]), .B1(p9_S[33]), .B2(
        p9_Partial_products_sum_add_23_n251), .C1(p9_C[32]), .C2(
        p9_Partial_products_sum_add_23_n251), .ZN(
        p9_Partial_products_sum_add_23_n248) );
  NAND2_X1 U3955 ( .A1(p9_Partial_products_sum_add_23_n252), .A2(
        p9_Partial_products_sum_add_23_n253), .ZN(
        p9_Partial_products_sum_add_23_n251) );
  OAI21_X1 U3956 ( .B1(p9_Partial_products_sum_add_23_n236), .B2(
        p9_Partial_products_sum_add_23_n237), .A(
        p9_Partial_products_sum_add_23_n238), .ZN(
        p9_Partial_products_sum_add_23_n235) );
  XNOR2_X1 U3957 ( .A(p9_Partial_products_sum_add_23_n196), .B(
        p9_Partial_products_sum_add_23_n199), .ZN(temp4[11]) );
  NOR2_X1 U3958 ( .A1(p9_C[41]), .A2(p9_S[42]), .ZN(
        p9_Partial_products_sum_add_23_n233) );
  NAND2_X1 U3959 ( .A1(p9_C[41]), .A2(p9_S[42]), .ZN(
        p9_Partial_products_sum_add_23_n234) );
  AOI222_X1 U3960 ( .A1(p9_Partial_products_sum_add_23_n235), .A2(p9_S[41]), 
        .B1(p9_Partial_products_sum_add_23_n235), .B2(p9_C[40]), .C1(p9_S[41]), 
        .C2(p9_C[40]), .ZN(p9_Partial_products_sum_add_23_n232) );
  XNOR2_X1 U3961 ( .A(p9_Partial_products_sum_add_23_n192), .B(
        p9_Partial_products_sum_add_23_n193), .ZN(temp4[13]) );
  NAND2_X1 U3962 ( .A1(p9_final_product2_25_), .A2(
        p9_Partial_products_sum_add_23_n194), .ZN(n3526) );
  AOI222_X1 U3963 ( .A1(p9_Partial_products_sum_add_23_n196), .A2(
        p9_Partial_products_sum_add_23_n197), .B1(
        p9_Partial_products_sum_add_23_n196), .B2(
        p9_Partial_products_sum_add_23_n198), .C1(
        p9_Partial_products_sum_add_23_n197), .C2(
        p9_Partial_products_sum_add_23_n198), .ZN(n3527) );
  AOI222_X1 U3964 ( .A1(p9_Partial_products_sum_add_23_n196), .A2(
        p9_Partial_products_sum_add_23_n197), .B1(
        p9_Partial_products_sum_add_23_n196), .B2(
        p9_Partial_products_sum_add_23_n198), .C1(
        p9_Partial_products_sum_add_23_n197), .C2(
        p9_Partial_products_sum_add_23_n198), .ZN(
        p9_Partial_products_sum_add_23_n194) );
  OAI21_X1 U3965 ( .B1(p9_Partial_products_sum_add_23_n203), .B2(
        p9_Partial_products_sum_add_23_n204), .A(
        p9_Partial_products_sum_add_23_n202), .ZN(n3530) );
  AOI222_X1 U3966 ( .A1(p9_Partial_products_sum_add_23_n208), .A2(
        p9_Partial_products_sum_add_23_n209), .B1(
        p9_Partial_products_sum_add_23_n208), .B2(
        p9_Partial_products_sum_add_23_n210), .C1(
        p9_Partial_products_sum_add_23_n209), .C2(
        p9_Partial_products_sum_add_23_n210), .ZN(
        p9_Partial_products_sum_add_23_n206) );
  OAI21_X1 U3967 ( .B1(p9_Partial_products_sum_add_23_n215), .B2(
        p9_Partial_products_sum_add_23_n216), .A(
        p9_Partial_products_sum_add_23_n214), .ZN(n3533) );
  AOI222_X1 U3968 ( .A1(p9_Partial_products_sum_add_23_n220), .A2(
        p9_Partial_products_sum_add_23_n221), .B1(
        p9_Partial_products_sum_add_23_n220), .B2(
        p9_Partial_products_sum_add_23_n222), .C1(
        p9_Partial_products_sum_add_23_n221), .C2(
        p9_Partial_products_sum_add_23_n222), .ZN(
        p9_Partial_products_sum_add_23_n218) );
  OAI21_X1 U3969 ( .B1(p9_Partial_products_sum_add_23_n227), .B2(
        p9_Partial_products_sum_add_23_n228), .A(
        p9_Partial_products_sum_add_23_n226), .ZN(n3536) );
  NAND2_X1 U3970 ( .A1(p9_Partial_products_sum_add_23_n230), .A2(p9_C[42]), 
        .ZN(n3537) );
  OAI21_X1 U3971 ( .B1(p9_Partial_products_sum_add_23_n230), .B2(p9_C[42]), 
        .A(p9_S[43]), .ZN(n3538) );
  NAND2_X1 U3972 ( .A1(p9_Partial_products_sum_add_23_n227), .A2(
        p9_Partial_products_sum_add_23_n228), .ZN(n3535) );
  AOI222_X1 U3973 ( .A1(p9_Partial_products_sum_add_23_n214), .A2(
        p9_Partial_products_sum_add_23_n215), .B1(
        p9_Partial_products_sum_add_23_n214), .B2(
        p9_Partial_products_sum_add_23_n216), .C1(
        p9_Partial_products_sum_add_23_n215), .C2(
        p9_Partial_products_sum_add_23_n216), .ZN(n3525) );
  NAND2_X1 U3974 ( .A1(p9_Partial_products_sum_add_23_n216), .A2(
        p9_Partial_products_sum_add_23_n215), .ZN(n3532) );
  NAND2_X1 U3975 ( .A1(p9_Partial_products_sum_add_23_n204), .A2(
        p9_Partial_products_sum_add_23_n203), .ZN(n3529) );
  AND2_X1 U3976 ( .A1(n3538), .A2(n3537), .ZN(
        p9_Partial_products_sum_add_23_n226) );
  AND2_X1 U3977 ( .A1(p9_S[45]), .A2(p9_C[44]), .ZN(n3541) );
  AND3_X1 U3978 ( .A1(n3536), .A2(p9_C[44]), .A3(n3535), .ZN(n3534) );
  AOI222_X1 U3979 ( .A1(p9_S[47]), .A2(p9_C[46]), .B1(p9_S[47]), .B2(n3521), 
        .C1(p9_C[46]), .C2(p9_Partial_products_sum_add_23_n218), .ZN(
        p9_Partial_products_sum_add_23_n214) );
  AND2_X1 U3980 ( .A1(p9_C[48]), .A2(p9_S[49]), .ZN(n3540) );
  AND3_X1 U3981 ( .A1(n3533), .A2(p9_C[48]), .A3(n3532), .ZN(n3531) );
  AND2_X1 U3982 ( .A1(p9_S[53]), .A2(p9_C[52]), .ZN(n3539) );
  AND3_X1 U3983 ( .A1(n3530), .A2(p9_C[52]), .A3(n3529), .ZN(n3528) );
  AOI222_X2 U3984 ( .A1(p9_Partial_products_sum_add_23_n202), .A2(
        p9_Partial_products_sum_add_23_n203), .B1(
        p9_Partial_products_sum_add_23_n202), .B2(
        p9_Partial_products_sum_add_23_n204), .C1(
        p9_Partial_products_sum_add_23_n203), .C2(
        p9_Partial_products_sum_add_23_n204), .ZN(n3522) );
  AOI211_X4 U3985 ( .C1(n3525), .C2(p9_S[49]), .A(n3540), .B(n3531), .ZN(
        p9_Partial_products_sum_add_23_n208) );
  AOI222_X2 U3986 ( .A1(p9_Partial_products_sum_add_23_n208), .A2(
        p9_Partial_products_sum_add_23_n209), .B1(
        p9_Partial_products_sum_add_23_n208), .B2(
        p9_Partial_products_sum_add_23_n210), .C1(
        p9_Partial_products_sum_add_23_n209), .C2(
        p9_Partial_products_sum_add_23_n210), .ZN(n3520) );
  AOI222_X4 U3987 ( .A1(p9_S[51]), .A2(p9_C[50]), .B1(n3520), .B2(p9_S[51]), 
        .C1(p9_C[50]), .C2(p9_Partial_products_sum_add_23_n206), .ZN(
        p9_Partial_products_sum_add_23_n202) );
  AOI222_X2 U3988 ( .A1(p9_Partial_products_sum_add_23_n226), .A2(
        p9_Partial_products_sum_add_23_n227), .B1(
        p9_Partial_products_sum_add_23_n226), .B2(
        p9_Partial_products_sum_add_23_n228), .C1(
        p9_Partial_products_sum_add_23_n227), .C2(
        p9_Partial_products_sum_add_23_n228), .ZN(n3519) );
  AOI211_X4 U3989 ( .C1(n3522), .C2(p9_S[53]), .A(n3539), .B(n3528), .ZN(
        p9_Partial_products_sum_add_23_n196) );
  NAND2_X1 U3990 ( .A1(p11_final_product1[1]), .A2(
        p11_Partial_products_sum_add_23_n318), .ZN(
        p11_Partial_products_sum_add_23_n315) );
  OAI21_X1 U3991 ( .B1(p11_Partial_products_sum_add_23_n307), .B2(
        p11_Partial_products_sum_add_23_n308), .A(
        p11_Partial_products_sum_add_23_n309), .ZN(
        p11_Partial_products_sum_add_23_n306) );
  OAI21_X1 U3992 ( .B1(p11_Partial_products_sum_add_23_n303), .B2(
        p11_Partial_products_sum_add_23_n304), .A(
        p11_Partial_products_sum_add_23_n305), .ZN(
        p11_Partial_products_sum_add_23_n302) );
  XNOR2_X1 U3993 ( .A(p11_Partial_products_sum_add_23_n276), .B(n3543), .ZN(
        temp6[6]) );
  XNOR2_X1 U3994 ( .A(p11_Partial_products_sum_add_23_n270), .B(
        p11_Partial_products_sum_add_23_n269), .ZN(temp6[8]) );
  XNOR2_X1 U3995 ( .A(p11_Partial_products_sum_add_23_n288), .B(
        p11_Partial_products_sum_add_23_n287), .ZN(temp6[2]) );
  XNOR2_X1 U3996 ( .A(p11_Partial_products_sum_add_23_n258), .B(n3545), .ZN(
        temp6[12]) );
  XNOR2_X1 U3997 ( .A(p11_Partial_products_sum_add_23_n264), .B(n3544), .ZN(
        temp6[10]) );
  AOI222_X1 U3998 ( .A1(p11_Partial_products_sum_add_23_n277), .A2(
        p11_Partial_products_sum_add_23_n278), .B1(
        p11_Partial_products_sum_add_23_n277), .B2(
        p11_Partial_products_sum_add_23_n279), .C1(
        p11_Partial_products_sum_add_23_n278), .C2(
        p11_Partial_products_sum_add_23_n279), .ZN(
        p11_Partial_products_sum_add_23_n275) );
  NOR2_X1 U3999 ( .A1(p11_C[37]), .A2(p11_S[38]), .ZN(
        p11_Partial_products_sum_add_23_n304) );
  AOI222_X1 U4000 ( .A1(p11_Partial_products_sum_add_23_n277), .A2(
        p11_Partial_products_sum_add_23_n278), .B1(
        p11_Partial_products_sum_add_23_n277), .B2(
        p11_Partial_products_sum_add_23_n279), .C1(
        p11_Partial_products_sum_add_23_n278), .C2(
        p11_Partial_products_sum_add_23_n279), .ZN(n3543) );
  NAND2_X1 U4001 ( .A1(p11_S[37]), .A2(p11_Partial_products_sum_add_23_n306), 
        .ZN(n3546) );
  NAND2_X1 U4002 ( .A1(p11_Partial_products_sum_add_23_n306), .A2(p11_C[36]), 
        .ZN(n3547) );
  NAND2_X1 U4003 ( .A1(p11_C[36]), .A2(p11_S[37]), .ZN(n3548) );
  AOI222_X1 U4004 ( .A1(p11_Partial_products_sum_add_23_n289), .A2(
        p11_Partial_products_sum_add_23_n290), .B1(
        p11_Partial_products_sum_add_23_n289), .B2(
        p11_Partial_products_sum_add_23_n291), .C1(
        p11_Partial_products_sum_add_23_n290), .C2(
        p11_Partial_products_sum_add_23_n291), .ZN(n3549) );
  OAI21_X1 U4005 ( .B1(p11_Partial_products_sum_add_23_n315), .B2(
        p11_Partial_products_sum_add_23_n316), .A(
        p11_Partial_products_sum_add_23_n317), .ZN(
        p11_Partial_products_sum_add_23_n314) );
  AOI222_X1 U4006 ( .A1(p11_S[33]), .A2(p11_C[32]), .B1(p11_S[33]), .B2(
        p11_Partial_products_sum_add_23_n314), .C1(p11_C[32]), .C2(
        p11_Partial_products_sum_add_23_n314), .ZN(
        p11_Partial_products_sum_add_23_n311) );
  OAI21_X1 U4007 ( .B1(p11_Partial_products_sum_add_23_n311), .B2(
        p11_Partial_products_sum_add_23_n312), .A(
        p11_Partial_products_sum_add_23_n313), .ZN(
        p11_Partial_products_sum_add_23_n310) );
  NAND2_X1 U4008 ( .A1(A1[3]), .A2(p11_S[32]), .ZN(
        p11_Partial_products_sum_add_23_n317) );
  NOR2_X1 U4009 ( .A1(A1[3]), .A2(p11_S[32]), .ZN(
        p11_Partial_products_sum_add_23_n316) );
  NAND2_X1 U4010 ( .A1(p11_C[34]), .A2(p11_Partial_products_sum_add_23_n310), 
        .ZN(n3550) );
  NAND2_X1 U4011 ( .A1(p11_S[35]), .A2(n3560), .ZN(n3551) );
  NAND2_X1 U4012 ( .A1(p11_S[35]), .A2(p11_C[34]), .ZN(n3552) );
  OAI21_X1 U4013 ( .B1(p11_Partial_products_sum_add_23_n299), .B2(
        p11_Partial_products_sum_add_23_n300), .A(
        p11_Partial_products_sum_add_23_n301), .ZN(
        p11_Partial_products_sum_add_23_n298) );
  NAND2_X1 U4014 ( .A1(p11_S[42]), .A2(p11_C[41]), .ZN(
        p11_Partial_products_sum_add_23_n297) );
  NOR2_X1 U4015 ( .A1(p11_S[42]), .A2(p11_C[41]), .ZN(
        p11_Partial_products_sum_add_23_n296) );
  NOR2_X1 U4016 ( .A1(p11_S[40]), .A2(p11_C[39]), .ZN(
        p11_Partial_products_sum_add_23_n300) );
  NAND2_X1 U4017 ( .A1(p11_S[40]), .A2(p11_C[39]), .ZN(
        p11_Partial_products_sum_add_23_n301) );
  NAND2_X1 U4018 ( .A1(p11_Partial_products_sum_add_23_n302), .A2(p11_C[38]), 
        .ZN(n3553) );
  NAND2_X1 U4019 ( .A1(p11_S[39]), .A2(p11_Partial_products_sum_add_23_n302), 
        .ZN(n3554) );
  NAND2_X1 U4020 ( .A1(p11_S[39]), .A2(p11_C[38]), .ZN(n3555) );
  XNOR2_X1 U4021 ( .A(p11_Partial_products_sum_add_23_n294), .B(n3559), .ZN(
        temp6[0]) );
  XNOR2_X1 U4022 ( .A(p11_Partial_products_sum_add_23_n277), .B(
        p11_Partial_products_sum_add_23_n280), .ZN(temp6[5]) );
  XNOR2_X1 U4023 ( .A(p11_Partial_products_sum_add_23_n283), .B(
        p11_Partial_products_sum_add_23_n286), .ZN(temp6[3]) );
  OAI21_X1 U4024 ( .B1(p11_Partial_products_sum_add_23_n296), .B2(
        p11_Partial_products_sum_add_23_n295), .A(
        p11_Partial_products_sum_add_23_n297), .ZN(
        p11_Partial_products_sum_add_23_n293) );
  NAND2_X1 U4025 ( .A1(p11_Partial_products_sum_add_23_n298), .A2(p11_C[40]), 
        .ZN(n3556) );
  NAND2_X1 U4026 ( .A1(p11_S[41]), .A2(n3561), .ZN(n3557) );
  NAND2_X1 U4027 ( .A1(p11_S[41]), .A2(p11_C[40]), .ZN(n3558) );
  XNOR2_X1 U4028 ( .A(p11_S[43]), .B(p11_C[42]), .ZN(
        p11_Partial_products_sum_add_23_n294) );
  NAND2_X1 U4029 ( .A1(p11_C[37]), .A2(p11_S[38]), .ZN(
        p11_Partial_products_sum_add_23_n305) );
  NOR2_X1 U4030 ( .A1(p11_C[33]), .A2(p11_S[34]), .ZN(
        p11_Partial_products_sum_add_23_n312) );
  XNOR2_X1 U4031 ( .A(p11_Partial_products_sum_add_23_n271), .B(
        p11_Partial_products_sum_add_23_n274), .ZN(temp6[7]) );
  XNOR2_X1 U4032 ( .A(p11_Partial_products_sum_add_23_n259), .B(
        p11_Partial_products_sum_add_23_n262), .ZN(temp6[11]) );
  XNOR2_X1 U4033 ( .A(p11_Partial_products_sum_add_23_n265), .B(
        p11_Partial_products_sum_add_23_n268), .ZN(temp6[9]) );
  XNOR2_X1 U4034 ( .A(p11_Partial_products_sum_add_23_n289), .B(
        p11_Partial_products_sum_add_23_n292), .ZN(temp6[1]) );
  NAND2_X1 U4035 ( .A1(p11_C[33]), .A2(p11_S[34]), .ZN(
        p11_Partial_products_sum_add_23_n313) );
  OAI21_X1 U4036 ( .B1(p11_Partial_products_sum_add_23_n311), .B2(
        p11_Partial_products_sum_add_23_n312), .A(
        p11_Partial_products_sum_add_23_n313), .ZN(n3560) );
  OAI21_X1 U4037 ( .B1(p11_Partial_products_sum_add_23_n299), .B2(
        p11_Partial_products_sum_add_23_n300), .A(
        p11_Partial_products_sum_add_23_n301), .ZN(n3561) );
  AOI22_X1 U4038 ( .A1(p11_S[44]), .A2(p11_C[43]), .B1(
        p11_Partial_products_sum_add_23_n291), .B2(
        p11_Partial_products_sum_add_23_n290), .ZN(
        p11_Partial_products_sum_add_23_n292) );
  NAND2_X1 U4039 ( .A1(n3564), .A2(n3563), .ZN(n3562) );
  XNOR2_X1 U4040 ( .A(n3570), .B(n3569), .ZN(temp6[13]) );
  NOR2_X1 U4041 ( .A1(n3562), .A2(p11_final_product2_26_), .ZN(n3567) );
  NOR2_X1 U4042 ( .A1(n3568), .A2(n3567), .ZN(n3570) );
  AOI21_X1 U4043 ( .B1(n3566), .B2(p11_final_product2_26_), .A(n3565), .ZN(
        n3568) );
  NAND2_X1 U4044 ( .A1(n3564), .A2(n3563), .ZN(n3566) );
  XOR2_X1 U4045 ( .A(p11_final_product2_26_), .B(p11_final_product1_26), .Z(
        n3569) );
  AOI222_X1 U4046 ( .A1(p11_Partial_products_sum_add_23_n265), .A2(
        p11_Partial_products_sum_add_23_n266), .B1(
        p11_Partial_products_sum_add_23_n265), .B2(
        p11_Partial_products_sum_add_23_n267), .C1(
        p11_Partial_products_sum_add_23_n266), .C2(
        p11_Partial_products_sum_add_23_n267), .ZN(
        p11_Partial_products_sum_add_23_n263) );
  NAND2_X1 U4047 ( .A1(n3572), .A2(n3571), .ZN(n3575) );
  OAI21_X1 U4048 ( .B1(p11_Partial_products_sum_add_23_n273), .B2(
        p11_Partial_products_sum_add_23_n272), .A(
        p11_Partial_products_sum_add_23_n271), .ZN(n3572) );
  NAND2_X1 U4049 ( .A1(p11_Partial_products_sum_add_23_n272), .A2(
        p11_Partial_products_sum_add_23_n273), .ZN(n3571) );
  NAND2_X1 U4050 ( .A1(p11_Partial_products_sum_add_23_n261), .A2(
        p11_Partial_products_sum_add_23_n260), .ZN(n3563) );
  AOI222_X1 U4051 ( .A1(p11_Partial_products_sum_add_23_n259), .A2(
        p11_Partial_products_sum_add_23_n260), .B1(
        p11_Partial_products_sum_add_23_n259), .B2(
        p11_Partial_products_sum_add_23_n261), .C1(
        p11_Partial_products_sum_add_23_n260), .C2(
        p11_Partial_products_sum_add_23_n261), .ZN(n3545) );
  AOI222_X1 U4052 ( .A1(p11_Partial_products_sum_add_23_n271), .A2(
        p11_Partial_products_sum_add_23_n272), .B1(
        p11_Partial_products_sum_add_23_n271), .B2(
        p11_Partial_products_sum_add_23_n273), .C1(
        p11_Partial_products_sum_add_23_n272), .C2(
        p11_Partial_products_sum_add_23_n273), .ZN(
        p11_Partial_products_sum_add_23_n269) );
  AND3_X1 U4053 ( .A1(n3552), .A2(n3551), .A3(n3550), .ZN(
        p11_Partial_products_sum_add_23_n307) );
  AND3_X1 U4054 ( .A1(n3548), .A2(n3547), .A3(n3546), .ZN(
        p11_Partial_products_sum_add_23_n303) );
  AND3_X1 U4055 ( .A1(n3558), .A2(n3557), .A3(n3556), .ZN(
        p11_Partial_products_sum_add_23_n295) );
  INV_X1 U4056 ( .A(p11_S[44]), .ZN(p11_Partial_products_sum_add_23_n290) );
  INV_X1 U4057 ( .A(p11_C[43]), .ZN(p11_Partial_products_sum_add_23_n291) );
  INV_X1 U4058 ( .A(p11_C[50]), .ZN(n3574) );
  INV_X1 U4059 ( .A(p11_S[51]), .ZN(n3573) );
  INV_X1 U4060 ( .A(p11_C[54]), .ZN(n3565) );
  AOI222_X4 U4061 ( .A1(p11_S[43]), .A2(p11_C[42]), .B1(n3559), .B2(p11_S[43]), 
        .C1(p11_Partial_products_sum_add_23_n293), .C2(p11_C[42]), .ZN(
        p11_Partial_products_sum_add_23_n289) );
  AOI222_X4 U4062 ( .A1(p11_S[45]), .A2(p11_C[44]), .B1(p11_S[45]), .B2(
        p11_Partial_products_sum_add_23_n287), .C1(p11_C[44]), .C2(n3549), 
        .ZN(p11_Partial_products_sum_add_23_n283) );
  AOI222_X4 U4063 ( .A1(p11_S[47]), .A2(p11_C[46]), .B1(p11_S[47]), .B2(
        p11_Partial_products_sum_add_23_n281), .C1(
        p11_Partial_products_sum_add_23_n281), .C2(p11_C[46]), .ZN(
        p11_Partial_products_sum_add_23_n277) );
  AOI222_X2 U4064 ( .A1(p11_Partial_products_sum_add_23_n289), .A2(
        p11_Partial_products_sum_add_23_n290), .B1(
        p11_Partial_products_sum_add_23_n289), .B2(
        p11_Partial_products_sum_add_23_n291), .C1(
        p11_Partial_products_sum_add_23_n290), .C2(
        p11_Partial_products_sum_add_23_n291), .ZN(
        p11_Partial_products_sum_add_23_n287) );
  AOI222_X1 U4065 ( .A1(p11_Partial_products_sum_add_23_n283), .A2(
        p11_Partial_products_sum_add_23_n284), .B1(
        p11_Partial_products_sum_add_23_n283), .B2(
        p11_Partial_products_sum_add_23_n285), .C1(
        p11_Partial_products_sum_add_23_n284), .C2(
        p11_Partial_products_sum_add_23_n285), .ZN(
        p11_Partial_products_sum_add_23_n281) );
  AOI222_X4 U4066 ( .A1(p11_S[49]), .A2(p11_C[48]), .B1(n3543), .B2(p11_S[49]), 
        .C1(p11_Partial_products_sum_add_23_n275), .C2(p11_C[48]), .ZN(
        p11_Partial_products_sum_add_23_n271) );
  AOI222_X1 U4067 ( .A1(p11_Partial_products_sum_add_23_n265), .A2(
        p11_Partial_products_sum_add_23_n266), .B1(
        p11_Partial_products_sum_add_23_n265), .B2(
        p11_Partial_products_sum_add_23_n267), .C1(
        p11_Partial_products_sum_add_23_n266), .C2(
        p11_Partial_products_sum_add_23_n267), .ZN(n3544) );
  AND3_X1 U4068 ( .A1(n3555), .A2(n3554), .A3(n3553), .ZN(
        p11_Partial_products_sum_add_23_n299) );
  AOI222_X4 U4069 ( .A1(p11_S[53]), .A2(p11_C[52]), .B1(n3544), .B2(p11_S[53]), 
        .C1(p11_Partial_products_sum_add_23_n263), .C2(p11_C[52]), .ZN(
        p11_Partial_products_sum_add_23_n259) );
  XNOR2_X1 U4070 ( .A(p10_Partial_products_sum_add_23_n306), .B(n3583), .ZN(
        temp5[4]) );
  XNOR2_X1 U4071 ( .A(p10_Partial_products_sum_add_23_n288), .B(
        p10_Partial_products_sum_add_23_n287), .ZN(temp5[10]) );
  XNOR2_X1 U4072 ( .A(p10_Partial_products_sum_add_23_n294), .B(n3577), .ZN(
        temp5[8]) );
  XNOR2_X1 U4073 ( .A(p10_Partial_products_sum_add_23_n312), .B(n3576), .ZN(
        temp5[2]) );
  OAI21_X1 U4074 ( .B1(p10_Partial_products_sum_add_23_n333), .B2(
        p10_Partial_products_sum_add_23_n334), .A(
        p10_Partial_products_sum_add_23_n335), .ZN(
        p10_Partial_products_sum_add_23_n332) );
  XNOR2_X1 U4075 ( .A(p10_Partial_products_sum_add_23_n300), .B(
        p10_Partial_products_sum_add_23_n299), .ZN(temp5[6]) );
  XNOR2_X1 U4076 ( .A(p10_Partial_products_sum_add_23_n313), .B(
        p10_Partial_products_sum_add_23_n316), .ZN(temp5[1]) );
  NAND2_X1 U4077 ( .A1(p10_Partial_products_sum_add_23_n327), .A2(
        p10_Partial_products_sum_add_23_n328), .ZN(
        p10_Partial_products_sum_add_23_n326) );
  OAI21_X1 U4078 ( .B1(p10_Partial_products_sum_add_23_n337), .B2(
        p10_Partial_products_sum_add_23_n338), .A(
        p10_Partial_products_sum_add_23_n339), .ZN(
        p10_Partial_products_sum_add_23_n336) );
  AOI222_X1 U4079 ( .A1(p10_Partial_products_sum_add_23_n313), .A2(
        p10_Partial_products_sum_add_23_n314), .B1(
        p10_Partial_products_sum_add_23_n313), .B2(
        p10_Partial_products_sum_add_23_n315), .C1(
        p10_Partial_products_sum_add_23_n314), .C2(
        p10_Partial_products_sum_add_23_n315), .ZN(n3576) );
  NAND2_X1 U4080 ( .A1(p10_C[38]), .A2(p10_Partial_products_sum_add_23_n326), 
        .ZN(n3578) );
  NAND2_X1 U4081 ( .A1(p10_S[39]), .A2(p10_Partial_products_sum_add_23_n326), 
        .ZN(n3579) );
  NAND2_X1 U4082 ( .A1(p10_C[34]), .A2(p10_Partial_products_sum_add_23_n336), 
        .ZN(n3580) );
  NAND2_X1 U4083 ( .A1(p10_Partial_products_sum_add_23_n336), .A2(p10_S[35]), 
        .ZN(n3581) );
  NAND2_X1 U4084 ( .A1(p10_S[35]), .A2(p10_C[34]), .ZN(n3582) );
  NOR2_X1 U4085 ( .A1(p10_C[33]), .A2(p10_S[34]), .ZN(
        p10_Partial_products_sum_add_23_n338) );
  XNOR2_X1 U4086 ( .A(p10_Partial_products_sum_add_23_n301), .B(
        p10_Partial_products_sum_add_23_n304), .ZN(temp5[5]) );
  NAND2_X1 U4087 ( .A1(p10_C[32]), .A2(p10_Partial_products_sum_add_23_n340), 
        .ZN(n3584) );
  NAND2_X1 U4088 ( .A1(p10_S[33]), .A2(p10_Partial_products_sum_add_23_n340), 
        .ZN(n3585) );
  NAND2_X1 U4089 ( .A1(p10_S[33]), .A2(p10_C[32]), .ZN(n3586) );
  XNOR2_X1 U4090 ( .A(p10_Partial_products_sum_add_23_n279), .B(
        p10_Partial_products_sum_add_23_n281), .ZN(temp5[12]) );
  XNOR2_X1 U4091 ( .A(p10_Partial_products_sum_add_23_n318), .B(
        p10_Partial_products_sum_add_23_n317), .ZN(temp5[0]) );
  NAND2_X1 U4092 ( .A1(p10_Partial_products_sum_add_23_n284), .A2(
        p10_Partial_products_sum_add_23_n285), .ZN(n3587) );
  NAND2_X1 U4093 ( .A1(p10_Partial_products_sum_add_23_n283), .A2(
        p10_Partial_products_sum_add_23_n285), .ZN(n3588) );
  NAND2_X1 U4094 ( .A1(p10_Partial_products_sum_add_23_n283), .A2(
        p10_Partial_products_sum_add_23_n284), .ZN(n3589) );
  XNOR2_X1 U4095 ( .A(p10_Partial_products_sum_add_23_n295), .B(
        p10_Partial_products_sum_add_23_n298), .ZN(temp5[7]) );
  XNOR2_X1 U4096 ( .A(n3597), .B(n3596), .ZN(temp5[13]) );
  NAND2_X1 U4097 ( .A1(n3594), .A2(n3595), .ZN(n3597) );
  OAI21_X1 U4098 ( .B1(p10_Partial_products_sum_add_23_n279), .B2(p10_C[54]), 
        .A(p10_final_product2_25_), .ZN(n3595) );
  NAND2_X1 U4099 ( .A1(p10_Partial_products_sum_add_23_n280), .A2(p10_C[53]), 
        .ZN(n3593) );
  NAND2_X1 U4100 ( .A1(p10_S[53]), .A2(p10_C[52]), .ZN(n3601) );
  NAND2_X1 U4101 ( .A1(p10_S[53]), .A2(n3598), .ZN(n3600) );
  NAND2_X1 U4102 ( .A1(p10_C[52]), .A2(n3602), .ZN(n3599) );
  AOI222_X1 U4103 ( .A1(p10_Partial_products_sum_add_23_n289), .A2(
        p10_Partial_products_sum_add_23_n290), .B1(
        p10_Partial_products_sum_add_23_n289), .B2(
        p10_Partial_products_sum_add_23_n291), .C1(
        p10_Partial_products_sum_add_23_n290), .C2(
        p10_Partial_products_sum_add_23_n291), .ZN(n3598) );
  AOI222_X1 U4104 ( .A1(p10_Partial_products_sum_add_23_n289), .A2(
        p10_Partial_products_sum_add_23_n290), .B1(
        p10_Partial_products_sum_add_23_n289), .B2(
        p10_Partial_products_sum_add_23_n291), .C1(
        p10_Partial_products_sum_add_23_n290), .C2(
        p10_Partial_products_sum_add_23_n291), .ZN(n3602) );
  OAI21_X1 U4105 ( .B1(p10_Partial_products_sum_add_23_n296), .B2(
        p10_Partial_products_sum_add_23_n297), .A(
        p10_Partial_products_sum_add_23_n295), .ZN(n3605) );
  NAND2_X1 U4106 ( .A1(p10_S[49]), .A2(p10_C[48]), .ZN(n3608) );
  NAND2_X1 U4107 ( .A1(p10_S[49]), .A2(p10_Partial_products_sum_add_23_n299), 
        .ZN(n3607) );
  NAND2_X1 U4108 ( .A1(p10_C[48]), .A2(n3609), .ZN(n3606) );
  AOI222_X1 U4109 ( .A1(p10_Partial_products_sum_add_23_n301), .A2(
        p10_Partial_products_sum_add_23_n302), .B1(
        p10_Partial_products_sum_add_23_n301), .B2(
        p10_Partial_products_sum_add_23_n303), .C1(
        p10_Partial_products_sum_add_23_n302), .C2(
        p10_Partial_products_sum_add_23_n303), .ZN(n3609) );
  OAI21_X1 U4110 ( .B1(p10_Partial_products_sum_add_23_n303), .B2(
        p10_Partial_products_sum_add_23_n302), .A(
        p10_Partial_products_sum_add_23_n301), .ZN(n3611) );
  NAND2_X1 U4111 ( .A1(p10_S[47]), .A2(p10_C[46]), .ZN(n3614) );
  NAND2_X1 U4112 ( .A1(p10_S[47]), .A2(n3615), .ZN(n3613) );
  NAND2_X1 U4113 ( .A1(p10_C[46]), .A2(p10_Partial_products_sum_add_23_n305), 
        .ZN(n3612) );
  AOI222_X1 U4114 ( .A1(p10_Partial_products_sum_add_23_n307), .A2(
        p10_Partial_products_sum_add_23_n308), .B1(
        p10_Partial_products_sum_add_23_n307), .B2(
        p10_Partial_products_sum_add_23_n309), .C1(
        p10_Partial_products_sum_add_23_n308), .C2(
        p10_Partial_products_sum_add_23_n309), .ZN(n3615) );
  AOI222_X1 U4115 ( .A1(p10_Partial_products_sum_add_23_n307), .A2(
        p10_Partial_products_sum_add_23_n308), .B1(
        p10_Partial_products_sum_add_23_n307), .B2(
        p10_Partial_products_sum_add_23_n309), .C1(
        p10_Partial_products_sum_add_23_n308), .C2(
        p10_Partial_products_sum_add_23_n309), .ZN(
        p10_Partial_products_sum_add_23_n305) );
  OAI21_X1 U4116 ( .B1(p10_Partial_products_sum_add_23_n314), .B2(
        p10_Partial_products_sum_add_23_n315), .A(
        p10_Partial_products_sum_add_23_n313), .ZN(n3618) );
  NAND2_X1 U4117 ( .A1(p10_Partial_products_sum_add_23_n317), .A2(p10_S[43]), 
        .ZN(n3620) );
  NAND2_X1 U4118 ( .A1(p10_Partial_products_sum_add_23_n317), .A2(p10_C[42]), 
        .ZN(n3621) );
  NAND2_X1 U4119 ( .A1(p10_S[43]), .A2(p10_C[42]), .ZN(n3619) );
  NAND2_X1 U4120 ( .A1(p10_Partial_products_sum_add_23_n314), .A2(
        p10_Partial_products_sum_add_23_n315), .ZN(n3617) );
  NAND2_X1 U4121 ( .A1(p10_Partial_products_sum_add_23_n303), .A2(
        p10_Partial_products_sum_add_23_n302), .ZN(n3610) );
  NAND2_X1 U4122 ( .A1(p10_Partial_products_sum_add_23_n296), .A2(
        p10_Partial_products_sum_add_23_n297), .ZN(n3622) );
  NAND2_X1 U4123 ( .A1(p10_Partial_products_sum_add_23_n296), .A2(
        p10_Partial_products_sum_add_23_n297), .ZN(n3604) );
  XNOR2_X1 U4124 ( .A(p10_final_product2_26_), .B(p10_final_product1_26), .ZN(
        n3596) );
  AOI222_X1 U4125 ( .A1(p10_Partial_products_sum_add_23_n289), .A2(
        p10_Partial_products_sum_add_23_n290), .B1(
        p10_Partial_products_sum_add_23_n289), .B2(
        p10_Partial_products_sum_add_23_n291), .C1(
        p10_Partial_products_sum_add_23_n290), .C2(
        p10_Partial_products_sum_add_23_n291), .ZN(
        p10_Partial_products_sum_add_23_n287) );
  AOI222_X1 U4126 ( .A1(p10_Partial_products_sum_add_23_n307), .A2(
        p10_Partial_products_sum_add_23_n308), .B1(
        p10_Partial_products_sum_add_23_n307), .B2(
        p10_Partial_products_sum_add_23_n309), .C1(
        p10_Partial_products_sum_add_23_n308), .C2(
        p10_Partial_products_sum_add_23_n309), .ZN(n3583) );
  INV_X1 U4127 ( .A(p10_S[48]), .ZN(p10_Partial_products_sum_add_23_n302) );
  AND2_X1 U4128 ( .A1(p10_S[41]), .A2(p10_C[40]), .ZN(n3592) );
  AND3_X1 U4129 ( .A1(n3586), .A2(n3585), .A3(n3584), .ZN(
        p10_Partial_products_sum_add_23_n337) );
  AND3_X1 U4130 ( .A1(n3582), .A2(n3581), .A3(n3580), .ZN(
        p10_Partial_products_sum_add_23_n333) );
  AND2_X1 U4131 ( .A1(p10_S[41]), .A2(p10_Partial_products_sum_add_23_n322), 
        .ZN(n3591) );
  AND2_X1 U4132 ( .A1(p10_C[40]), .A2(p10_Partial_products_sum_add_23_n322), 
        .ZN(n3590) );
  AND2_X1 U4133 ( .A1(p10_S[45]), .A2(p10_C[44]), .ZN(n3624) );
  AND3_X1 U4134 ( .A1(n3618), .A2(p10_C[44]), .A3(n3617), .ZN(n3616) );
  AND2_X1 U4135 ( .A1(n3611), .A2(n3610), .ZN(
        p10_Partial_products_sum_add_23_n299) );
  AND2_X1 U4136 ( .A1(p10_C[50]), .A2(p10_S[51]), .ZN(n3625) );
  AND3_X1 U4137 ( .A1(n3605), .A2(p10_C[50]), .A3(n3604), .ZN(n3603) );
  INV_X1 U4138 ( .A(p10_Partial_products_sum_add_23_n283), .ZN(
        p10_Partial_products_sum_add_23_n280) );
  INV_X1 U4139 ( .A(p10_C[53]), .ZN(p10_Partial_products_sum_add_23_n284) );
  INV_X1 U4140 ( .A(p10_S[54]), .ZN(p10_Partial_products_sum_add_23_n285) );
  AND3_X1 U4141 ( .A1(n3589), .A2(n3588), .A3(n3587), .ZN(
        p10_Partial_products_sum_add_23_n279) );
  INV_X1 U4142 ( .A(p10_C[54]), .ZN(p10_Partial_products_sum_add_23_n277) );
  AOI211_X4 U4143 ( .C1(n3576), .C2(p10_S[45]), .A(n3624), .B(n3616), .ZN(
        p10_Partial_products_sum_add_23_n307) );
  AOI211_X4 U4144 ( .C1(n3577), .C2(p10_S[51]), .A(n3625), .B(n3603), .ZN(
        p10_Partial_products_sum_add_23_n289) );
  AND3_X2 U4145 ( .A1(n3614), .A2(n3613), .A3(n3612), .ZN(
        p10_Partial_products_sum_add_23_n301) );
  AND2_X2 U4146 ( .A1(n3623), .A2(n3622), .ZN(n3577) );
  NAND2_X1 U4147 ( .A1(n3626), .A2(p10_Partial_products_sum_add_23_n295), .ZN(
        n3623) );
  OR2_X1 U4148 ( .A1(p10_Partial_products_sum_add_23_n297), .A2(
        p10_Partial_products_sum_add_23_n296), .ZN(n3626) );
  AND3_X2 U4149 ( .A1(n3621), .A2(n3620), .A3(n3619), .ZN(
        p10_Partial_products_sum_add_23_n313) );
  AOI222_X1 U4150 ( .A1(p6_Partial_products_sum_add_23_n194), .A2(
        p6_Partial_products_sum_add_23_n195), .B1(
        p6_Partial_products_sum_add_23_n194), .B2(
        p6_Partial_products_sum_add_23_n196), .C1(
        p6_Partial_products_sum_add_23_n195), .C2(
        p6_Partial_products_sum_add_23_n196), .ZN(
        p6_Partial_products_sum_add_23_n192) );
  OAI21_X1 U4151 ( .B1(p6_Partial_products_sum_add_23_n228), .B2(
        p6_Partial_products_sum_add_23_n229), .A(
        p6_Partial_products_sum_add_23_n230), .ZN(
        p6_Partial_products_sum_add_23_n227) );
  OAI21_X1 U4152 ( .B1(p6_Partial_products_sum_add_23_n224), .B2(
        p6_Partial_products_sum_add_23_n225), .A(
        p6_Partial_products_sum_add_23_n226), .ZN(
        p6_Partial_products_sum_add_23_n223) );
  OAI21_X1 U4153 ( .B1(p6_Partial_products_sum_add_23_n220), .B2(
        p6_Partial_products_sum_add_23_n221), .A(
        p6_Partial_products_sum_add_23_n222), .ZN(
        p6_Partial_products_sum_add_23_n219) );
  XNOR2_X1 U4154 ( .A(p6_Partial_products_sum_add_23_n193), .B(n3627), .ZN(
        temp1[6]) );
  XNOR2_X1 U4155 ( .A(p6_Partial_products_sum_add_23_n174), .B(
        p6_Partial_products_sum_add_23_n175), .ZN(temp1[12]) );
  NAND2_X1 U4156 ( .A1(p6_S[35]), .A2(p6_C[34]), .ZN(n3628) );
  NAND2_X1 U4157 ( .A1(p6_Partial_products_sum_add_23_n227), .A2(p6_C[34]), 
        .ZN(n3629) );
  NAND2_X1 U4158 ( .A1(p6_Partial_products_sum_add_23_n227), .A2(p6_S[35]), 
        .ZN(n3630) );
  NAND2_X1 U4159 ( .A1(p6_S[37]), .A2(p6_C[36]), .ZN(n3631) );
  NAND2_X1 U4160 ( .A1(p6_Partial_products_sum_add_23_n223), .A2(p6_C[36]), 
        .ZN(n3632) );
  NAND2_X1 U4161 ( .A1(p6_Partial_products_sum_add_23_n223), .A2(p6_S[37]), 
        .ZN(n3633) );
  XNOR2_X1 U4162 ( .A(n3641), .B(p6_Partial_products_sum_add_23_n203), .ZN(
        temp1[3]) );
  XNOR2_X1 U4163 ( .A(p6_Partial_products_sum_add_23_n181), .B(n3635), .ZN(
        temp1[10]) );
  XNOR2_X1 U4164 ( .A(p6_Partial_products_sum_add_23_n187), .B(n3636), .ZN(
        temp1[8]) );
  XNOR2_X1 U4165 ( .A(p6_Partial_products_sum_add_23_n199), .B(n3634), .ZN(
        temp1[4]) );
  OAI21_X1 U4166 ( .B1(p6_Partial_products_sum_add_23_n216), .B2(
        p6_Partial_products_sum_add_23_n217), .A(
        p6_Partial_products_sum_add_23_n218), .ZN(
        p6_Partial_products_sum_add_23_n215) );
  AOI222_X1 U4167 ( .A1(p6_Partial_products_sum_add_23_n219), .A2(p6_S[39]), 
        .B1(p6_Partial_products_sum_add_23_n219), .B2(p6_C[38]), .C1(p6_S[39]), 
        .C2(p6_C[38]), .ZN(p6_Partial_products_sum_add_23_n216) );
  AOI222_X1 U4168 ( .A1(n3640), .A2(p6_Partial_products_sum_add_23_n201), .B1(
        n3640), .B2(p6_Partial_products_sum_add_23_n202), .C1(
        p6_Partial_products_sum_add_23_n201), .C2(
        p6_Partial_products_sum_add_23_n202), .ZN(
        p6_Partial_products_sum_add_23_n198) );
  NAND2_X1 U4169 ( .A1(p6_Partial_products_sum_add_23_n232), .A2(
        p6_Partial_products_sum_add_23_n233), .ZN(
        p6_Partial_products_sum_add_23_n231) );
  AOI222_X1 U4170 ( .A1(p6_S[33]), .A2(p6_C[32]), .B1(p6_S[33]), .B2(
        p6_Partial_products_sum_add_23_n231), .C1(p6_C[32]), .C2(
        p6_Partial_products_sum_add_23_n231), .ZN(
        p6_Partial_products_sum_add_23_n228) );
  AOI222_X1 U4171 ( .A1(n3641), .A2(p6_Partial_products_sum_add_23_n201), .B1(
        p6_Partial_products_sum_add_23_n200), .B2(
        p6_Partial_products_sum_add_23_n202), .C1(
        p6_Partial_products_sum_add_23_n201), .C2(
        p6_Partial_products_sum_add_23_n202), .ZN(n3634) );
  XNOR2_X1 U4172 ( .A(p6_Partial_products_sum_add_23_n188), .B(
        p6_Partial_products_sum_add_23_n191), .ZN(temp1[7]) );
  AOI222_X1 U4173 ( .A1(p6_S[45]), .A2(p6_C[44]), .B1(p6_S[45]), .B2(
        p6_Partial_products_sum_add_23_n204), .C1(p6_C[44]), .C2(
        p6_Partial_products_sum_add_23_n204), .ZN(
        p6_Partial_products_sum_add_23_n200) );
  NAND2_X1 U4174 ( .A1(p6_S[41]), .A2(p6_C[40]), .ZN(n3637) );
  NAND2_X1 U4175 ( .A1(p6_Partial_products_sum_add_23_n215), .A2(p6_C[40]), 
        .ZN(n3638) );
  NAND2_X1 U4176 ( .A1(p6_Partial_products_sum_add_23_n215), .A2(p6_S[41]), 
        .ZN(n3639) );
  AOI222_X1 U4177 ( .A1(p6_S[45]), .A2(p6_C[44]), .B1(p6_S[45]), .B2(
        p6_Partial_products_sum_add_23_n204), .C1(p6_C[44]), .C2(
        p6_Partial_products_sum_add_23_n204), .ZN(n3641) );
  AOI222_X1 U4178 ( .A1(p6_S[45]), .A2(p6_C[44]), .B1(p6_S[45]), .B2(
        p6_Partial_products_sum_add_23_n204), .C1(p6_C[44]), .C2(
        p6_Partial_products_sum_add_23_n204), .ZN(n3640) );
  XNOR2_X1 U4179 ( .A(n3642), .B(n3643), .ZN(temp1[13]) );
  XOR2_X1 U4180 ( .A(p6_final_product2_26_), .B(p6_final_product1_26), .Z(
        n3643) );
  NAND2_X1 U4181 ( .A1(p6_Partial_products_sum_add_23_n174), .A2(p6_C[54]), 
        .ZN(n3645) );
  NAND2_X1 U4182 ( .A1(p6_Partial_products_sum_add_23_n174), .A2(
        p6_final_product2_25_), .ZN(n3646) );
  AOI222_X1 U4183 ( .A1(p6_Partial_products_sum_add_23_n182), .A2(
        p6_Partial_products_sum_add_23_n183), .B1(
        p6_Partial_products_sum_add_23_n182), .B2(
        p6_Partial_products_sum_add_23_n184), .C1(
        p6_Partial_products_sum_add_23_n183), .C2(
        p6_Partial_products_sum_add_23_n184), .ZN(
        p6_Partial_products_sum_add_23_n180) );
  AOI21_X1 U4184 ( .B1(n3651), .B2(n3650), .A(n3649), .ZN(n3653) );
  NAND2_X1 U4185 ( .A1(n3648), .A2(n3647), .ZN(n3651) );
  OAI21_X1 U4186 ( .B1(p6_Partial_products_sum_add_23_n190), .B2(
        p6_Partial_products_sum_add_23_n189), .A(
        p6_Partial_products_sum_add_23_n188), .ZN(n3648) );
  NAND2_X1 U4187 ( .A1(p6_Partial_products_sum_add_23_n189), .A2(
        p6_Partial_products_sum_add_23_n190), .ZN(n3647) );
  NAND2_X1 U4188 ( .A1(p6_C[54]), .A2(p6_final_product2_25_), .ZN(n3644) );
  AOI222_X1 U4189 ( .A1(p6_Partial_products_sum_add_23_n188), .A2(
        p6_Partial_products_sum_add_23_n189), .B1(
        p6_Partial_products_sum_add_23_n188), .B2(
        p6_Partial_products_sum_add_23_n190), .C1(
        p6_Partial_products_sum_add_23_n189), .C2(
        p6_Partial_products_sum_add_23_n190), .ZN(n3636) );
  NOR2_X1 U4190 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  AND3_X1 U4191 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(
        p6_Partial_products_sum_add_23_n224) );
  AND3_X1 U4192 ( .A1(n3633), .A2(n3632), .A3(n3631), .ZN(
        p6_Partial_products_sum_add_23_n220) );
  INV_X1 U4193 ( .A(p6_C[50]), .ZN(n3650) );
  INV_X1 U4194 ( .A(p6_S[51]), .ZN(n3649) );
  NOR2_X1 U4195 ( .A1(n3653), .A2(n3652), .ZN(
        p6_Partial_products_sum_add_23_n182) );
  AND3_X1 U4196 ( .A1(n3645), .A2(n3646), .A3(n3644), .ZN(n3642) );
  AOI222_X4 U4197 ( .A1(p6_S[43]), .A2(p6_C[42]), .B1(p6_S[43]), .B2(
        p6_Partial_products_sum_add_23_n210), .C1(p6_C[42]), .C2(
        p6_Partial_products_sum_add_23_n210), .ZN(
        p6_Partial_products_sum_add_23_n206) );
  AOI222_X2 U4198 ( .A1(p6_Partial_products_sum_add_23_n206), .A2(
        p6_Partial_products_sum_add_23_n207), .B1(
        p6_Partial_products_sum_add_23_n206), .B2(
        p6_Partial_products_sum_add_23_n208), .C1(
        p6_Partial_products_sum_add_23_n207), .C2(
        p6_Partial_products_sum_add_23_n208), .ZN(
        p6_Partial_products_sum_add_23_n204) );
  AOI222_X4 U4199 ( .A1(p6_S[49]), .A2(p6_C[48]), .B1(p6_S[49]), .B2(n3627), 
        .C1(p6_Partial_products_sum_add_23_n192), .C2(p6_C[48]), .ZN(
        p6_Partial_products_sum_add_23_n188) );
  AOI222_X4 U4200 ( .A1(p6_S[47]), .A2(p6_C[46]), .B1(p6_S[47]), .B2(n3634), 
        .C1(p6_C[46]), .C2(p6_Partial_products_sum_add_23_n198), .ZN(
        p6_Partial_products_sum_add_23_n194) );
  AOI222_X2 U4201 ( .A1(p6_Partial_products_sum_add_23_n176), .A2(
        p6_Partial_products_sum_add_23_n177), .B1(
        p6_Partial_products_sum_add_23_n176), .B2(
        p6_Partial_products_sum_add_23_n178), .C1(
        p6_Partial_products_sum_add_23_n177), .C2(
        p6_Partial_products_sum_add_23_n178), .ZN(
        p6_Partial_products_sum_add_23_n174) );
  AOI222_X1 U4202 ( .A1(p6_Partial_products_sum_add_23_n182), .A2(
        p6_Partial_products_sum_add_23_n183), .B1(
        p6_Partial_products_sum_add_23_n182), .B2(
        p6_Partial_products_sum_add_23_n184), .C1(
        p6_Partial_products_sum_add_23_n183), .C2(
        p6_Partial_products_sum_add_23_n184), .ZN(n3635) );
  AOI222_X2 U4203 ( .A1(p6_Partial_products_sum_add_23_n194), .A2(
        p6_Partial_products_sum_add_23_n195), .B1(
        p6_Partial_products_sum_add_23_n194), .B2(
        p6_Partial_products_sum_add_23_n196), .C1(
        p6_Partial_products_sum_add_23_n195), .C2(
        p6_Partial_products_sum_add_23_n196), .ZN(n3627) );
  AND3_X2 U4204 ( .A1(n3657), .A2(n3656), .A3(n3655), .ZN(
        p6_Partial_products_sum_add_23_n176) );
  NAND2_X1 U4205 ( .A1(p6_S[53]), .A2(n3635), .ZN(n3656) );
  NAND2_X1 U4206 ( .A1(p6_S[53]), .A2(p6_C[52]), .ZN(n3657) );
  INV_X2 U4207 ( .A(B3[10]), .ZN(n642) );
  XOR2_X1 U4208 ( .A(n2387), .B(n2390), .Z(n3658) );
  XOR2_X1 U4209 ( .A(n3825), .B(n3658), .Z(p11_S[42]) );
  INV_X2 U4210 ( .A(B3[5]), .ZN(n714) );
  NAND2_X1 U4211 ( .A1(n3659), .A2(n2472), .ZN(n2757) );
  AOI211_X4 U4212 ( .C1(reg3_reg[5]), .C2(reg3_reg[6]), .A(n3696), .B(n1404), 
        .ZN(n1149) );
  AOI221_X1 U4213 ( .B1(n1884), .B2(B0[10]), .C1(n1885), .C2(n1991), .A(n2237), 
        .ZN(n2236) );
  NAND2_X2 U4214 ( .A1(n3803), .A2(A1[3]), .ZN(n2561) );
  XNOR2_X1 U4215 ( .A(n2716), .B(n3660), .ZN(n2713) );
  XOR2_X1 U4216 ( .A(n2714), .B(n2711), .Z(n3660) );
  AOI211_X4 U4217 ( .C1(A2[7]), .C2(A2[8]), .A(n3158), .B(n3179), .ZN(n2907)
         );
  INV_X2 U4218 ( .A(B2[10]), .ZN(n1092) );
  INV_X1 U4219 ( .A(n2472), .ZN(n3661) );
  INV_X2 U4220 ( .A(n3661), .ZN(n3662) );
  INV_X2 U4221 ( .A(B2[5]), .ZN(n1164) );
  AOI211_X4 U4222 ( .C1(reg1_reg[1]), .C2(reg1_reg[2]), .A(n3717), .B(n2322), 
        .ZN(n2149) );
  XNOR2_X1 U4223 ( .A(n3663), .B(n2675), .ZN(n2676) );
  XOR2_X1 U4224 ( .A(n2678), .B(n2679), .Z(n3663) );
  AOI211_X4 U4225 ( .C1(reg2_reg[1]), .C2(reg2_reg[2]), .A(n3718), .B(n1872), 
        .ZN(n1699) );
  AOI211_X4 U4226 ( .C1(A2[7]), .C2(A2[8]), .A(A2[9]), .B(n3179), .ZN(n2906)
         );
  AOI211_X4 U4227 ( .C1(A1[7]), .C2(A1[8]), .A(n2712), .B(n2733), .ZN(n2457)
         );
  AOI211_X4 U4228 ( .C1(A2[3]), .C2(A2[4]), .A(A2[5]), .B(n3212), .ZN(n2984)
         );
  AOI211_X4 U4229 ( .C1(A2[4]), .C2(A2[3]), .A(n2873), .B(n3212), .ZN(n2985)
         );
  AOI211_X4 U4230 ( .C1(A2[6]), .C2(A2[5]), .A(A2[7]), .B(n3203), .ZN(n2947)
         );
  AOI211_X4 U4231 ( .C1(A1[3]), .C2(A1[4]), .A(A1[5]), .B(n2766), .ZN(n2531)
         );
  AOI211_X4 U4232 ( .C1(reg3_reg[1]), .C2(reg3_reg[2]), .A(reg3_reg[3]), .B(
        n1422), .ZN(n1249) );
  AOI211_X4 U4233 ( .C1(A1[4]), .C2(A1[3]), .A(n2423), .B(n2766), .ZN(n2532)
         );
  AOI211_X4 U4234 ( .C1(A2[1]), .C2(A2[2]), .A(n3213), .B(n3219), .ZN(n3048)
         );
  AOI211_X4 U4235 ( .C1(A2[1]), .C2(A2[2]), .A(A2[3]), .B(n3219), .ZN(n3047)
         );
  AOI211_X4 U4236 ( .C1(reg4_reg[1]), .C2(reg4_reg[2]), .A(n3703), .B(n973), 
        .ZN(n800) );
  NAND2_X2 U4237 ( .A1(A1[7]), .A2(A1[8]), .ZN(n2447) );
  AOI211_X4 U4238 ( .C1(A1[7]), .C2(A1[8]), .A(A1[9]), .B(n2733), .ZN(n2456)
         );
  AOI211_X4 U4239 ( .C1(A1[6]), .C2(A1[5]), .A(A1[7]), .B(n2757), .ZN(n2497)
         );
  NAND2_X2 U4240 ( .A1(A2[6]), .A2(A2[5]), .ZN(n2922) );
  AOI211_X4 U4241 ( .C1(A2[5]), .C2(A2[6]), .A(n2859), .B(n3203), .ZN(n2948)
         );
  AOI211_X4 U4242 ( .C1(A1[5]), .C2(A1[6]), .A(n2409), .B(n2757), .ZN(n2498)
         );
  INV_X1 U4243 ( .A(VIN), .ZN(n3849) );
  INV_X1 U4244 ( .A(VIN), .ZN(n3850) );
  INV_X1 U4245 ( .A(VIN), .ZN(n3846) );
  INV_X1 U4246 ( .A(VIN), .ZN(n3851) );
  INV_X1 U4247 ( .A(VIN), .ZN(n3847) );
  INV_X1 U4248 ( .A(n2832), .ZN(n3821) );
  AND2_X1 U4249 ( .A1(n2948), .A2(n3678), .ZN(n3843) );
  AND2_X1 U4250 ( .A1(n2947), .A2(reg4[6]), .ZN(n3842) );
  INV_X1 U4251 ( .A(n2840), .ZN(n3822) );
  INV_X1 U4252 ( .A(n2921), .ZN(n3202) );
  AND2_X1 U4253 ( .A1(A2[3]), .A2(n3219), .ZN(n3709) );
  INV_X1 U4254 ( .A(n3159), .ZN(n3176) );
  INV_X1 U4255 ( .A(n2896), .ZN(n3178) );
  NAND2_X1 U4256 ( .A1(n3203), .A2(A2[7]), .ZN(n2921) );
  INV_X1 U4257 ( .A(A2[11]), .ZN(n3120) );
  NAND2_X1 U4258 ( .A1(A2[9]), .A2(A2[10]), .ZN(n2880) );
  NAND2_X1 U4259 ( .A1(A2[11]), .A2(A2[12]), .ZN(n2776) );
  INV_X1 U4260 ( .A(VIN), .ZN(n3852) );
  INV_X1 U4261 ( .A(p6_final_product2_26_), .ZN(p6_final_product2_25_) );
  INV_X1 U4262 ( .A(n1932), .ZN(n3820) );
  INV_X1 U4263 ( .A(n2226), .ZN(n3780) );
  AND2_X1 U4264 ( .A1(B0[7]), .A2(n2148), .ZN(n3784) );
  AND2_X1 U4265 ( .A1(B0[2]), .A2(n2112), .ZN(n3779) );
  AND2_X1 U4266 ( .A1(B0[3]), .A2(n2148), .ZN(n3726) );
  AND2_X1 U4267 ( .A1(n1969), .A2(n1970), .ZN(n3809) );
  INV_X1 U4268 ( .A(n1882), .ZN(n3777) );
  AND2_X1 U4269 ( .A1(B0[2]), .A2(n1884), .ZN(n3794) );
  INV_X1 U4270 ( .A(n2111), .ZN(n3783) );
  AND2_X1 U4271 ( .A1(B0[0]), .A2(n2148), .ZN(n3786) );
  INV_X1 U4272 ( .A(n2195), .ZN(n2205) );
  INV_X1 U4273 ( .A(n2194), .ZN(n3824) );
  OR2_X1 U4274 ( .A1(n2003), .A2(n2112), .ZN(n3832) );
  INV_X1 U4275 ( .A(n2131), .ZN(n2128) );
  INV_X1 U4276 ( .A(n2139), .ZN(n2136) );
  INV_X1 U4277 ( .A(n1889), .ZN(n1884) );
  INV_X1 U4278 ( .A(p8_final_product2_26_), .ZN(p8_final_product2_25_) );
  INV_X1 U4279 ( .A(n1045), .ZN(n3811) );
  INV_X1 U4280 ( .A(n1048), .ZN(n3805) );
  INV_X1 U4281 ( .A(n1374), .ZN(n1054) );
  INV_X1 U4282 ( .A(n983), .ZN(n3816) );
  OR2_X1 U4283 ( .A1(n3787), .A2(n3788), .ZN(n3791) );
  INV_X1 U4284 ( .A(n1232), .ZN(n1229) );
  INV_X1 U4285 ( .A(n1254), .ZN(n1253) );
  INV_X1 U4286 ( .A(n1240), .ZN(n1237) );
  INV_X1 U4287 ( .A(n990), .ZN(n985) );
  INV_X1 U4288 ( .A(n782), .ZN(n779) );
  NOR2_X1 U4289 ( .A1(n783), .A2(n582), .ZN(n578) );
  INV_X1 U4290 ( .A(n583), .ZN(n3810) );
  INV_X1 U4291 ( .A(n845), .ZN(n3813) );
  INV_X1 U4292 ( .A(n592), .ZN(n3806) );
  INV_X1 U4293 ( .A(n877), .ZN(n3799) );
  OR2_X1 U4294 ( .A1(n692), .A2(n763), .ZN(n3831) );
  OR2_X1 U4295 ( .A1(B3[6]), .A2(n762), .ZN(n3830) );
  INV_X1 U4296 ( .A(n603), .ZN(n3815) );
  INV_X1 U4297 ( .A(n533), .ZN(n3812) );
  INV_X1 U4298 ( .A(n790), .ZN(n787) );
  INV_X1 U4299 ( .A(n540), .ZN(n535) );
  INV_X1 U4300 ( .A(p9_final_product2_26_), .ZN(p9_final_product2_25_) );
  INV_X1 U4301 ( .A(VIN), .ZN(n3848) );
  INV_X1 U4302 ( .A(n1482), .ZN(n3800) );
  INV_X1 U4303 ( .A(n1494), .ZN(n3814) );
  INV_X1 U4304 ( .A(n1776), .ZN(n3798) );
  INV_X1 U4305 ( .A(n1824), .ZN(n1503) );
  INV_X1 U4306 ( .A(n1849), .ZN(n1514) );
  INV_X1 U4307 ( .A(n1527), .ZN(n3795) );
  CLKBUF_X1 U4308 ( .A(n1489), .Z(n3829) );
  INV_X1 U4309 ( .A(n1744), .ZN(n3797) );
  INV_X1 U4310 ( .A(n1742), .ZN(n3785) );
  INV_X1 U4311 ( .A(n1681), .ZN(n1678) );
  NOR2_X1 U4312 ( .A1(n1682), .A2(n1481), .ZN(n1477) );
  INV_X1 U4313 ( .A(n1439), .ZN(n1434) );
  INV_X1 U4314 ( .A(p7_final_product2_26_), .ZN(p7_final_product2_25_) );
  INV_X1 U4315 ( .A(p11_final_product2_26_), .ZN(p11_final_product2_25_) );
  INV_X1 U4316 ( .A(n2382), .ZN(n3808) );
  AND2_X1 U4317 ( .A1(n2742), .A2(n2743), .ZN(n2741) );
  INV_X1 U4318 ( .A(n2561), .ZN(n2747) );
  INV_X1 U4319 ( .A(n2713), .ZN(n2730) );
  INV_X1 U4320 ( .A(n2446), .ZN(n2732) );
  INV_X1 U4321 ( .A(n2676), .ZN(n2695) );
  OR2_X1 U4322 ( .A1(n3687), .A2(n2562), .ZN(n3835) );
  OR2_X1 U4323 ( .A1(reg2[6]), .A2(n2561), .ZN(n3834) );
  AND2_X1 U4324 ( .A1(n3844), .A2(n3845), .ZN(n3828) );
  OR2_X1 U4325 ( .A1(n2648), .A2(n2444), .ZN(n3844) );
  OR2_X1 U4326 ( .A1(reg2[9]), .A2(n2561), .ZN(n3838) );
  OR2_X1 U4327 ( .A1(n3691), .A2(n2562), .ZN(n3839) );
  INV_X1 U4328 ( .A(n2581), .ZN(n2578) );
  XOR2_X1 U4329 ( .A(n2610), .B(n2583), .Z(n2381) );
  INV_X1 U4330 ( .A(n2590), .ZN(n2587) );
  INV_X1 U4331 ( .A(A1[5]), .ZN(n2423) );
  CLKBUF_X1 U4332 ( .A(n2518), .Z(n3826) );
  OAI21_X1 U4333 ( .B1(A1[3]), .B2(A1[4]), .A(n2518), .ZN(n2766) );
  NAND2_X1 U4334 ( .A1(A1[9]), .A2(A1[10]), .ZN(n2430) );
  INV_X1 U4335 ( .A(A1[13]), .ZN(n2444) );
  NAND2_X1 U4336 ( .A1(A1[11]), .A2(A1[12]), .ZN(n2326) );
  NOR2_X1 U4337 ( .A1(n2132), .A2(n1931), .ZN(n1927) );
  NAND2_X1 U4338 ( .A1(A1[1]), .A2(A1[2]), .ZN(n2562) );
  NAND2_X1 U4339 ( .A1(A2[3]), .A2(A2[4]), .ZN(n2968) );
  NAND2_X1 U4340 ( .A1(A2[1]), .A2(A2[2]), .ZN(n3009) );
  NAND2_X1 U4341 ( .A1(A1[1]), .A2(n2771), .ZN(n2332) );
  AOI222_X1 U4342 ( .A1(n3840), .A2(n2840), .B1(n3840), .B2(n2837), .C1(n2840), 
        .C2(n2837), .ZN(p10_C[42]) );
  NAND2_X1 U4343 ( .A1(n3118), .A2(n3117), .ZN(n3817) );
  NAND2_X1 U4344 ( .A1(n2864), .A2(n2863), .ZN(n3819) );
  AOI222_X1 U4345 ( .A1(n2847), .A2(n2848), .B1(n2847), .B2(n2845), .C1(n2848), 
        .C2(n2845), .ZN(p10_C[40]) );
  XOR2_X1 U4346 ( .A(n3142), .B(n3121), .Z(n3122) );
  NAND2_X1 U4347 ( .A1(A2[1]), .A2(n3218), .ZN(n2782) );
  AOI222_X1 U4348 ( .A1(n2823), .A2(n2824), .B1(n2823), .B2(n2821), .C1(n2824), 
        .C2(n2821), .ZN(p10_C[46]) );
  AOI222_X1 U4349 ( .A1(n2815), .A2(n2816), .B1(n2815), .B2(n2813), .C1(n2816), 
        .C2(n2813), .ZN(p10_C[48]) );
  AOI222_X1 U4350 ( .A1(n2892), .A2(n2893), .B1(n2892), .B2(n2798), .C1(n2893), 
        .C2(n2798), .ZN(p10_C[52]) );
  AOI222_X1 U4351 ( .A1(n1951), .A2(n1952), .B1(n1951), .B2(n1949), .C1(n1952), 
        .C2(n1949), .ZN(p6_C[39]) );
  NAND2_X1 U4352 ( .A1(n2005), .A2(n3777), .ZN(n3776) );
  NAND2_X1 U4353 ( .A1(B0[9]), .A2(n1884), .ZN(n3775) );
  NAND2_X1 U4354 ( .A1(n2041), .A2(n3783), .ZN(n3782) );
  AOI221_X1 U4355 ( .B1(n2148), .B2(B0[5]), .C1(n2149), .C2(n2063), .A(n2297), 
        .ZN(n2275) );
  AOI222_X1 U4356 ( .A1(n1974), .A2(n3711), .B1(n1974), .B2(n1972), .C1(n3711), 
        .C2(n1972), .ZN(p6_C[34]) );
  AOI211_X1 U4357 ( .C1(n2133), .C2(n1885), .A(n3794), .B(n3793), .ZN(n1978)
         );
  AOI211_X1 U4358 ( .C1(n1888), .C2(n2149), .A(n3786), .B(n3783), .ZN(n1977)
         );
  AOI222_X1 U4359 ( .A1(n3833), .A2(n1940), .B1(n3833), .B2(n1937), .C1(n1940), 
        .C2(n1937), .ZN(p6_C[42]) );
  AOI221_X1 U4360 ( .B1(n2047), .B2(B0[5]), .C1(n2048), .C2(n2063), .A(n2231), 
        .ZN(n2203) );
  AOI221_X1 U4361 ( .B1(n2148), .B2(B0[9]), .C1(n2149), .C2(n2003), .A(n2242), 
        .ZN(n2219) );
  AOI221_X1 U4362 ( .B1(n2047), .B2(B0[9]), .C1(n2048), .C2(n2003), .A(n2145), 
        .ZN(n2104) );
  AOI222_X1 U4363 ( .A1(n1044), .A2(n1045), .B1(n1044), .B2(n1042), .C1(n1045), 
        .C2(n1042), .ZN(p8_C[41]) );
  XNOR2_X1 U4364 ( .A(n1049), .B(n3805), .ZN(n3804) );
  AOI222_X1 U4365 ( .A1(n1052), .A2(n1053), .B1(n1052), .B2(n1050), .C1(n1053), 
        .C2(n1050), .ZN(p8_C[39]) );
  AOI221_X1 U4366 ( .B1(n1249), .B2(B2[5]), .C1(n1250), .C2(n1164), .A(n1397), 
        .ZN(n1375) );
  AOI222_X1 U4367 ( .A1(n1075), .A2(n3698), .B1(n1075), .B2(n1073), .C1(n3698), 
        .C2(n1073), .ZN(p8_C[34]) );
  AOI221_X1 U4368 ( .B1(n986), .B2(n1092), .C1(n985), .C2(B2[10]), .A(n1337), 
        .ZN(n1336) );
  AOI221_X1 U4369 ( .B1(B2[8]), .B2(n1249), .C1(n1250), .C2(n1106), .A(n1338), 
        .ZN(n1335) );
  AOI221_X1 U4370 ( .B1(n1148), .B2(B2[5]), .C1(n1149), .C2(n1164), .A(n1331), 
        .ZN(n1304) );
  AOI221_X1 U4371 ( .B1(n1249), .B2(B2[9]), .C1(n1250), .C2(n1104), .A(n1342), 
        .ZN(n1318) );
  NAND2_X1 U4372 ( .A1(B2[10]), .A2(n1249), .ZN(n3790) );
  OAI221_X1 U4373 ( .B1(B2[2]), .B2(n975), .C1(n1234), .C2(n977), .A(n1235), 
        .ZN(n1222) );
  AOI222_X1 U4374 ( .A1(n582), .A2(n583), .B1(n582), .B2(n580), .C1(n583), 
        .C2(n580), .ZN(p9_C[44]) );
  AOI222_X1 U4375 ( .A1(n590), .A2(n591), .B1(n590), .B2(n588), .C1(n591), 
        .C2(n588), .ZN(p9_C[42]) );
  AOI222_X1 U4376 ( .A1(n870), .A2(n871), .B1(n871), .B2(n872), .C1(n870), 
        .C2(n872), .ZN(n862) );
  AOI222_X1 U4377 ( .A1(n594), .A2(n595), .B1(n594), .B2(n592), .C1(n595), 
        .C2(n592), .ZN(p9_C[41]) );
  AOI221_X1 U4378 ( .B1(n536), .B2(n642), .C1(n535), .C2(B3[10]), .A(n888), 
        .ZN(n887) );
  AOI222_X1 U4379 ( .A1(n602), .A2(n603), .B1(n602), .B2(n600), .C1(n603), 
        .C2(n600), .ZN(p9_C[39]) );
  AOI221_X1 U4380 ( .B1(n799), .B2(B3[5]), .C1(n800), .C2(n714), .A(n948), 
        .ZN(n926) );
  AOI222_X1 U4381 ( .A1(n625), .A2(n3699), .B1(n625), .B2(n623), .C1(n3699), 
        .C2(n623), .ZN(p9_C[34]) );
  AOI221_X1 U4382 ( .B1(n698), .B2(B3[9]), .C1(n699), .C2(n654), .A(n796), 
        .ZN(n755) );
  AOI222_X1 U4383 ( .A1(n543), .A2(n544), .B1(n543), .B2(n542), .C1(n544), 
        .C2(n542), .ZN(p9_C[54]) );
  AOI221_X1 U4384 ( .B1(n1698), .B2(B1[5]), .C1(n1699), .C2(n1613), .A(n1847), 
        .ZN(n1825) );
  AOI222_X1 U4385 ( .A1(n1524), .A2(n3712), .B1(n1524), .B2(n1522), .C1(n3712), 
        .C2(n1522), .ZN(p7_C[34]) );
  AOI222_X1 U4386 ( .A1(n3829), .A2(n1490), .B1(n3829), .B2(n1487), .C1(n1490), 
        .C2(n1487), .ZN(p7_C[42]) );
  AOI221_X1 U4387 ( .B1(n1597), .B2(B1[5]), .C1(n1598), .C2(n1613), .A(n1781), 
        .ZN(n1753) );
  AOI222_X1 U4388 ( .A1(n1769), .A2(n1770), .B1(n1770), .B2(n1771), .C1(n1769), 
        .C2(n1771), .ZN(n1761) );
  AOI222_X1 U4389 ( .A1(n1481), .A2(n1482), .B1(n1481), .B2(n1479), .C1(n1482), 
        .C2(n1479), .ZN(p7_C[44]) );
  AOI222_X1 U4390 ( .A1(n1465), .A2(n1466), .B1(n1465), .B2(n1463), .C1(n1466), 
        .C2(n1463), .ZN(p7_C[48]) );
  AOI222_X1 U4391 ( .A1(n1442), .A2(n1443), .B1(n1442), .B2(n1441), .C1(n1443), 
        .C2(n1441), .ZN(p7_C[54]) );
  AOI222_X1 U4392 ( .A1(n2342), .A2(n2343), .B1(n2342), .B2(n2341), .C1(n2343), 
        .C2(n2341), .ZN(p11_C[54]) );
  AOI222_X1 U4393 ( .A1(n2424), .A2(n2423), .B1(n2424), .B2(n2422), .C1(n2423), 
        .C2(n2422), .ZN(p11_C[34]) );
  AOI221_X1 U4394 ( .B1(n2456), .B2(reg2[0]), .C1(n2457), .C2(n3689), .A(n2732), .ZN(n2711) );
  AOI222_X1 U4395 ( .A1(n3828), .A2(n2390), .B1(n3828), .B2(n2387), .C1(n2390), 
        .C2(n2387), .ZN(p11_C[42]) );
  AOI221_X1 U4396 ( .B1(n2531), .B2(reg2[7]), .C1(n2532), .C2(n3688), .A(n2692), .ZN(n2672) );
  NAND3_X1 U4397 ( .A1(n3774), .A2(n3775), .A3(n3776), .ZN(n2250) );
  NAND2_X1 U4398 ( .A1(n2003), .A2(n1885), .ZN(n3774) );
  AOI21_X1 U4399 ( .B1(n2133), .B2(n2111), .A(n3779), .ZN(n3778) );
  AOI211_X1 U4400 ( .C1(n2149), .C2(n2115), .A(n3726), .B(n3778), .ZN(n2299)
         );
  FA_X1 U4401 ( .A(n2223), .B(n3780), .CI(n2227), .S(n2224) );
  XNOR2_X1 U4402 ( .A(n1504), .B(n1824), .ZN(p7_S[38]) );
  AOI21_X1 U4403 ( .B1(n2017), .B2(n2149), .A(n3784), .ZN(n3781) );
  OAI211_X1 U4404 ( .C1(n2041), .C2(n2112), .A(n3781), .B(n3782), .ZN(n2251)
         );
  XNOR2_X1 U4405 ( .A(n2251), .B(n2250), .ZN(n2256) );
  XNOR2_X1 U4406 ( .A(n1743), .B(n3785), .ZN(n1747) );
  OAI22_X1 U4407 ( .A1(n1104), .A2(n1213), .B1(B2[9]), .B2(n1212), .ZN(n3787)
         );
  NAND2_X1 U4408 ( .A1(n1092), .A2(n1250), .ZN(n3789) );
  NAND2_X1 U4409 ( .A1(n3789), .A2(n3790), .ZN(n3788) );
  XNOR2_X1 U4410 ( .A(n3791), .B(n1281), .ZN(n1283) );
  XNOR2_X1 U4411 ( .A(n1283), .B(n1292), .ZN(n1312) );
  XNOR2_X1 U4412 ( .A(n1312), .B(n1282), .ZN(n1294) );
  XNOR2_X1 U4413 ( .A(n2182), .B(n2191), .ZN(n3792) );
  XNOR2_X1 U4414 ( .A(n3792), .B(n2181), .ZN(n2193) );
  NOR2_X1 U4415 ( .A1(B0[1]), .A2(n1882), .ZN(n3793) );
  XNOR2_X1 U4416 ( .A(n1528), .B(n3795), .ZN(p7_S[32]) );
  FA_X1 U4417 ( .A(n2199), .B(n2203), .CI(n2204), .S(n2201) );
  XNOR2_X1 U4418 ( .A(n1941), .B(n1942), .ZN(p6_S[41]) );
  XNOR2_X1 U4419 ( .A(n833), .B(n842), .ZN(n3796) );
  XNOR2_X1 U4420 ( .A(n3796), .B(n832), .ZN(n844) );
  FA_X1 U4421 ( .A(n904), .B(n908), .CI(n909), .S(n906) );
  XOR2_X1 U4422 ( .A(n605), .B(n604), .Z(p9_S[38]) );
  FA_X1 U4423 ( .A(n1746), .B(n3797), .CI(n1748), .S(n1745) );
  FA_X1 U4424 ( .A(n1773), .B(n3798), .CI(n1777), .S(n1774) );
  FA_X1 U4425 ( .A(n1803), .B(n1807), .CI(n1808), .S(n1805) );
  XNOR2_X1 U4426 ( .A(n1499), .B(n1500), .ZN(p7_S[39]) );
  FA_X1 U4427 ( .A(n874), .B(n3799), .CI(n878), .S(n875) );
  XNOR2_X1 U4428 ( .A(n1487), .B(n1488), .ZN(p7_S[42]) );
  FA_X1 U4429 ( .A(n1479), .B(n3800), .CI(n1481), .S(p7_S[44]) );
  XOR2_X1 U4430 ( .A(n2262), .B(n2259), .Z(n3801) );
  XNOR2_X1 U4431 ( .A(n2264), .B(n3801), .ZN(n2261) );
  XNOR2_X1 U4432 ( .A(n1949), .B(n1950), .ZN(p6_S[39]) );
  OAI22_X1 U4433 ( .A1(n2332), .A2(reg2[1]), .B1(reg2[2]), .B2(n2337), .ZN(
        n3802) );
  AOI21_X1 U4434 ( .B1(n2334), .B2(reg2[2]), .A(n3802), .ZN(n2427) );
  XNOR2_X1 U4435 ( .A(A1[1]), .B(A1[2]), .ZN(n3803) );
  XNOR2_X1 U4436 ( .A(n2659), .B(n2649), .ZN(n2648) );
  AOI222_X1 U4437 ( .A1(n2219), .A2(n2220), .B1(n2220), .B2(n2221), .C1(n2219), 
        .C2(n2221), .ZN(n2211) );
  XNOR2_X1 U4438 ( .A(n1046), .B(n3804), .ZN(p8_S[40]) );
  XNOR2_X1 U4439 ( .A(n594), .B(n595), .ZN(n3807) );
  XNOR2_X1 U4440 ( .A(n3807), .B(n3806), .ZN(p9_S[41]) );
  FA_X1 U4441 ( .A(n2379), .B(n3808), .CI(n2381), .S(p11_S[44]) );
  FA_X1 U4442 ( .A(n1965), .B(n3809), .CI(n1967), .S(p6_S[35]) );
  FA_X1 U4443 ( .A(n580), .B(n3810), .CI(n582), .S(p9_S[44]) );
  FA_X1 U4444 ( .A(n1042), .B(n3811), .CI(n1044), .S(p8_S[41]) );
  XNOR2_X1 U4445 ( .A(A2[1]), .B(A2[2]), .ZN(n3219) );
  XNOR2_X1 U4446 ( .A(n1945), .B(n1946), .ZN(p6_S[40]) );
  AOI221_X1 U4447 ( .B1(n3689), .B2(n2602), .C1(reg2[0]), .C2(n2601), .A(n2747), .ZN(n2428) );
  FA_X1 U4448 ( .A(n847), .B(n3813), .CI(n849), .S(n846) );
  FA_X1 U4449 ( .A(n1491), .B(n3814), .CI(n1493), .S(p7_S[41]) );
  FA_X1 U4450 ( .A(n600), .B(n3815), .CI(n602), .S(p9_S[39]) );
  XNOR2_X1 U4451 ( .A(n1495), .B(n1496), .ZN(p7_S[40]) );
  XOR2_X1 U4452 ( .A(n2428), .B(n2427), .Z(p11_S[32]) );
  AOI221_X1 U4453 ( .B1(n2947), .B2(reg4[0]), .C1(n2948), .C2(n3670), .A(n3202), .ZN(n3188) );
  XNOR2_X1 U4454 ( .A(n3188), .B(n3189), .ZN(n2861) );
  XOR2_X1 U4455 ( .A(n1307), .B(n1297), .Z(n3818) );
  AOI22_X1 U4456 ( .A1(n1296), .A2(n3761), .B1(n3818), .B2(reg3_reg[13]), .ZN(
        n1040) );
  XNOR2_X1 U4457 ( .A(n1038), .B(n1039), .ZN(p8_S[42]) );
  FA_X1 U4458 ( .A(n1353), .B(n1357), .CI(n1358), .S(n1355) );
  XNOR2_X1 U4459 ( .A(n1050), .B(n1051), .ZN(p8_S[39]) );
  FA_X1 U4460 ( .A(n2859), .B(n3819), .CI(n2861), .S(p10_S[36]) );
  XOR2_X1 U4461 ( .A(n3105), .B(n3095), .Z(n3841) );
  FA_X1 U4462 ( .A(n3151), .B(n3155), .CI(n3156), .S(n3153) );
  XNOR2_X1 U4463 ( .A(n2845), .B(n2846), .ZN(p10_S[40]) );
  XNOR2_X1 U4464 ( .A(n1055), .B(n1374), .ZN(p8_S[38]) );
  XNOR2_X1 U4465 ( .A(n596), .B(n597), .ZN(p9_S[40]) );
  FA_X1 U4466 ( .A(n1929), .B(n3820), .CI(n1931), .S(p6_S[44]) );
  XNOR2_X1 U4467 ( .A(n589), .B(n588), .ZN(p9_S[42]) );
  FA_X1 U4468 ( .A(n2829), .B(n3821), .CI(n2831), .S(p10_S[44]) );
  FA_X1 U4469 ( .A(n2837), .B(n3822), .CI(n3823), .S(p10_S[42]) );
  AOI22_X1 U4470 ( .A1(n3094), .A2(n2894), .B1(n3841), .B2(A2[13]), .ZN(n3823)
         );
  FA_X1 U4471 ( .A(n2196), .B(n3824), .CI(n2198), .S(n2195) );
  AOI22_X1 U4472 ( .A1(reg1_reg[13]), .A2(n2205), .B1(n2195), .B2(n3757), .ZN(
        n1939) );
  XNOR2_X1 U4473 ( .A(n1937), .B(n1938), .ZN(p6_S[42]) );
  NAND2_X1 U4474 ( .A1(n3844), .A2(n3845), .ZN(n3825) );
  XNOR2_X1 U4475 ( .A(n3240), .B(reg7[13]), .ZN(SUB1_N13) );
  XNOR2_X1 U4476 ( .A(n2867), .B(n2868), .ZN(n2866) );
  NAND2_X1 U4477 ( .A1(n2867), .A2(n2865), .ZN(n3205) );
  OAI211_X1 U4478 ( .C1(n2867), .C2(n2865), .A(n2870), .B(n2869), .ZN(n3204)
         );
  XOR2_X1 U4479 ( .A(n2864), .B(n2863), .Z(n2867) );
  AOI22_X1 U4480 ( .A1(reg4[2]), .A2(n3047), .B1(n3048), .B2(n3673), .ZN(n3209) );
  AOI22_X1 U4481 ( .A1(n787), .A2(n788), .B1(n789), .B2(n790), .ZN(n777) );
  XNOR2_X1 U4482 ( .A(n3110), .B(n3081), .ZN(n3092) );
  OAI221_X1 U4483 ( .B1(reg2[13]), .B2(n2446), .C1(n3680), .C2(n2447), .A(
        n2448), .ZN(n2445) );
  OAI221_X1 U4484 ( .B1(reg2[12]), .B2(n2446), .C1(n3690), .C2(n2447), .A(
        n2448), .ZN(n2349) );
  AOI22_X1 U4485 ( .A1(reg2[11]), .A2(n2447), .B1(n2446), .B2(n3686), .ZN(
        n2474) );
  AOI22_X1 U4486 ( .A1(reg2[10]), .A2(n2447), .B1(n2446), .B2(n3693), .ZN(
        n2496) );
  OAI221_X1 U4487 ( .B1(reg2[8]), .B2(n2446), .C1(n3683), .C2(n2447), .A(n2530), .ZN(n2529) );
  AOI22_X1 U4488 ( .A1(reg2[9]), .A2(n2447), .B1(n2446), .B2(n3691), .ZN(n2516) );
  OAI221_X1 U4489 ( .B1(reg2[5]), .B2(n2446), .C1(n3677), .C2(n2447), .A(n2620), .ZN(n2589) );
  AOI22_X1 U4490 ( .A1(reg2[0]), .A2(n2447), .B1(n2446), .B2(n3689), .ZN(n2717) );
  AOI22_X1 U4491 ( .A1(reg2[2]), .A2(n2447), .B1(n2446), .B2(n3692), .ZN(n2682) );
  AOI22_X1 U4492 ( .A1(reg2[4]), .A2(n2447), .B1(n2446), .B2(n3685), .ZN(n2637) );
  AOI22_X1 U4493 ( .A1(reg2[7]), .A2(n2447), .B1(n2446), .B2(n3688), .ZN(n2564) );
  AOI22_X1 U4494 ( .A1(reg2[1]), .A2(n2447), .B1(n2446), .B2(n3684), .ZN(n2704) );
  AOI22_X1 U4495 ( .A1(reg2[6]), .A2(n2447), .B1(n2446), .B2(n3687), .ZN(n2599) );
  AOI22_X1 U4496 ( .A1(reg2[3]), .A2(n2447), .B1(n2446), .B2(n3669), .ZN(n2663) );
  NAND2_X1 U4497 ( .A1(A1[3]), .A2(A1[4]), .ZN(n2518) );
  OAI211_X1 U4498 ( .C1(A2[7]), .C2(n2861), .A(n2864), .B(n2863), .ZN(n3199)
         );
  AOI22_X1 U4499 ( .A1(reg2[13]), .A2(n2531), .B1(n2532), .B2(n3680), .ZN(
        n2519) );
  AOI22_X1 U4500 ( .A1(reg2[12]), .A2(n2531), .B1(n2532), .B2(n3690), .ZN(
        n2560) );
  AOI221_X1 U4501 ( .B1(n2531), .B2(reg2[11]), .C1(n2532), .C2(n3686), .A(
        n2603), .ZN(n2600) );
  AOI221_X1 U4502 ( .B1(n2531), .B2(reg2[10]), .C1(n2532), .C2(n3693), .A(
        n2622), .ZN(n2593) );
  AOI221_X1 U4503 ( .B1(n2531), .B2(reg2[5]), .C1(n2532), .C2(n3677), .A(n2724), .ZN(n2709) );
  AOI221_X1 U4504 ( .B1(n2531), .B2(reg2[4]), .C1(n2532), .C2(n3685), .A(n2738), .ZN(n2735) );
  AOI221_X1 U4505 ( .B1(n2531), .B2(reg2[2]), .C1(n2532), .C2(n3692), .A(n2755), .ZN(n2743) );
  AOI22_X1 U4506 ( .A1(reg2[1]), .A2(n2531), .B1(n2532), .B2(n3684), .ZN(n2760) );
  XNOR2_X1 U4507 ( .A(n2470), .B(n2464), .ZN(n2465) );
  AOI22_X1 U4508 ( .A1(n2459), .A2(n2460), .B1(n2461), .B2(n2462), .ZN(n2354)
         );
  OAI21_X1 U4509 ( .B1(n2534), .B2(n2535), .A(n2536), .ZN(n2528) );
  OAI211_X1 U4510 ( .C1(n618), .C2(n616), .A(n621), .B(n620), .ZN(n956) );
  NAND2_X1 U4511 ( .A1(n618), .A2(n616), .ZN(n957) );
  AOI22_X1 U4512 ( .A1(reg4[7]), .A2(n3047), .B1(n3048), .B2(n3672), .ZN(n3167) );
  AOI22_X1 U4513 ( .A1(A1[11]), .A2(n2676), .B1(n2695), .B2(n2674), .ZN(n2395)
         );
  AOI22_X1 U4514 ( .A1(reg2[13]), .A2(n2497), .B1(n2498), .B2(n3680), .ZN(
        n2473) );
  AOI22_X1 U4515 ( .A1(reg2[10]), .A2(n2497), .B1(n2498), .B2(n3693), .ZN(
        n2558) );
  AOI221_X1 U4516 ( .B1(n2497), .B2(reg2[2]), .C1(n2498), .C2(n3692), .A(n2734), .ZN(n2714) );
  AOI221_X1 U4517 ( .B1(n2497), .B2(reg2[0]), .C1(n2498), .C2(n3689), .A(n2756), .ZN(n2742) );
  AOI222_X1 U4518 ( .A1(n1048), .A2(n1049), .B1(n1048), .B2(n1046), .C1(n1049), 
        .C2(n1046), .ZN(p8_C[40]) );
  XNOR2_X1 U4519 ( .A(n2608), .B(n2609), .ZN(n2631) );
  NAND2_X1 U4520 ( .A1(n2616), .A2(n2618), .ZN(n2617) );
  XNOR2_X1 U4521 ( .A(n2616), .B(n2618), .ZN(n2638) );
  OAI22_X1 U4522 ( .A1(n1252), .A2(n1253), .B1(n1254), .B2(n1255), .ZN(n1243)
         );
  AOI22_X1 U4523 ( .A1(B2[10]), .A2(n977), .B1(n975), .B2(n1092), .ZN(n1091)
         );
  AOI22_X1 U4524 ( .A1(B2[10]), .A2(n1081), .B1(n1080), .B2(n1092), .ZN(n1109)
         );
  AOI221_X1 U4525 ( .B1(n1089), .B2(B2[10]), .C1(n1090), .C2(n1092), .A(n1120), 
        .ZN(n1114) );
  AOI22_X1 U4526 ( .A1(B2[10]), .A2(n1098), .B1(n1097), .B2(n1092), .ZN(n1147)
         );
  AOI221_X1 U4527 ( .B1(n1107), .B2(B2[10]), .C1(n1108), .C2(n1092), .A(n1167), 
        .ZN(n1153) );
  AOI22_X1 U4528 ( .A1(B2[10]), .A2(n1123), .B1(n1122), .B2(n1092), .ZN(n1184)
         );
  AOI22_X1 U4529 ( .A1(B2[10]), .A2(n1148), .B1(n1149), .B2(n1092), .ZN(n1209)
         );
  NAND2_X1 U4530 ( .A1(A1[7]), .A2(n2411), .ZN(n2754) );
  OAI211_X1 U4531 ( .C1(A1[7]), .C2(n2411), .A(n2414), .B(n2413), .ZN(n2753)
         );
  XNOR2_X1 U4532 ( .A(n2411), .B(n2412), .ZN(n2410) );
  AOI222_X1 U4533 ( .A1(n1947), .A2(n1948), .B1(n1947), .B2(n1945), .C1(n1948), 
        .C2(n1945), .ZN(p6_C[40]) );
  NAND3_X1 U4534 ( .A1(n3830), .A2(n3831), .A3(n920), .ZN(n902) );
  AOI221_X1 U4535 ( .B1(n1148), .B2(B2[2]), .C1(n1149), .C2(n1234), .A(n1382), 
        .ZN(n1362) );
  OAI221_X1 U4536 ( .B1(B1[6]), .B2(n1661), .C1(n1591), .C2(n1662), .A(n1819), 
        .ZN(n1801) );
  XNOR2_X1 U4537 ( .A(n1801), .B(n1800), .ZN(n1806) );
  AOI22_X1 U4538 ( .A1(B3[6]), .A2(n799), .B1(n800), .B2(n692), .ZN(n936) );
  AOI22_X1 U4539 ( .A1(B3[6]), .A2(n719), .B1(n718), .B2(n692), .ZN(n891) );
  AOI221_X1 U4540 ( .B1(n698), .B2(B3[6]), .C1(n699), .C2(n692), .A(n866), 
        .ZN(n842) );
  XNOR2_X1 U4541 ( .A(n2742), .B(n2743), .ZN(n2411) );
  AOI22_X1 U4542 ( .A1(n884), .A2(n885), .B1(n886), .B2(n887), .ZN(n883) );
  AOI222_X1 U4543 ( .A1(n598), .A2(n599), .B1(n598), .B2(n596), .C1(n599), 
        .C2(n596), .ZN(p9_C[40]) );
  AOI22_X1 U4544 ( .A1(reg2[2]), .A2(n2601), .B1(n2602), .B2(n3692), .ZN(n2763) );
  AOI22_X1 U4545 ( .A1(reg2[3]), .A2(n2601), .B1(n2602), .B2(n3669), .ZN(n2762) );
  AOI22_X1 U4546 ( .A1(reg2[6]), .A2(n2601), .B1(n2602), .B2(n3687), .ZN(n2737) );
  AOI22_X1 U4547 ( .A1(n2587), .A2(n2588), .B1(n2589), .B2(n2590), .ZN(n2576)
         );
  NAND2_X1 U4548 ( .A1(n1350), .A2(n1351), .ZN(n1347) );
  AOI22_X1 U4549 ( .A1(n1678), .A2(n1679), .B1(n1680), .B2(n1681), .ZN(n1476)
         );
  AOI22_X1 U4550 ( .A1(n779), .A2(n780), .B1(n781), .B2(n782), .ZN(n577) );
  XNOR2_X1 U4551 ( .A(n812), .B(n783), .ZN(n582) );
  AOI22_X1 U4552 ( .A1(reg1_reg[13]), .A2(n2205), .B1(n2195), .B2(n3757), .ZN(
        n3833) );
  AOI22_X1 U4553 ( .A1(n2136), .A2(n2137), .B1(n2138), .B2(n2139), .ZN(n2126)
         );
  NAND3_X1 U4554 ( .A1(n3834), .A2(n3835), .A3(n2721), .ZN(n2703) );
  XNOR2_X1 U4555 ( .A(n2391), .B(n2392), .ZN(p11_S[41]) );
  AOI22_X1 U4556 ( .A1(B2[8]), .A2(n977), .B1(n975), .B2(n1106), .ZN(n1105) );
  AOI22_X1 U4557 ( .A1(B2[8]), .A2(n979), .B1(n980), .B2(n1106), .ZN(n1119) );
  AOI22_X1 U4558 ( .A1(B2[8]), .A2(n1081), .B1(n1080), .B2(n1106), .ZN(n1146)
         );
  AOI221_X1 U4559 ( .B1(n1089), .B2(B2[8]), .C1(n1090), .C2(n1106), .A(n1165), 
        .ZN(n1140) );
  OAI221_X1 U4560 ( .B1(B2[8]), .B2(n1097), .C1(n1106), .C2(n1098), .A(n1181), 
        .ZN(n1180) );
  AOI221_X1 U4561 ( .B1(n1107), .B2(B2[8]), .C1(n1108), .C2(n1106), .A(n1215), 
        .ZN(n1190) );
  AOI22_X1 U4562 ( .A1(B2[8]), .A2(n1123), .B1(n1122), .B2(n1106), .ZN(n1246)
         );
  OAI221_X1 U4563 ( .B1(B2[8]), .B2(n1168), .C1(n1106), .C2(n1169), .A(n1286), 
        .ZN(n1276) );
  AOI22_X1 U4564 ( .A1(B2[8]), .A2(n1213), .B1(n1212), .B2(n1106), .ZN(n1342)
         );
  AOI22_X1 U4565 ( .A1(B2[8]), .A2(n985), .B1(n986), .B2(n1106), .ZN(n1384) );
  XNOR2_X1 U4566 ( .A(n2664), .B(n2635), .ZN(n2646) );
  NAND2_X1 U4567 ( .A1(n901), .A2(n902), .ZN(n898) );
  XNOR2_X1 U4568 ( .A(n902), .B(n901), .ZN(n907) );
  XNOR2_X1 U4569 ( .A(n1326), .B(n1327), .ZN(n1344) );
  AOI221_X1 U4570 ( .B1(n979), .B2(B2[5]), .C1(n980), .C2(n1164), .A(n1175), 
        .ZN(n1154) );
  AOI22_X1 U4571 ( .A1(B2[5]), .A2(n977), .B1(n975), .B2(n1164), .ZN(n1163) );
  OAI221_X1 U4572 ( .B1(B2[5]), .B2(n1080), .C1(n1164), .C2(n1081), .A(n1207), 
        .ZN(n1193) );
  OAI221_X1 U4573 ( .B1(B2[5]), .B2(n1097), .C1(n1164), .C2(n1098), .A(n1267), 
        .ZN(n1239) );
  AOI22_X1 U4574 ( .A1(B2[5]), .A2(n1107), .B1(n1108), .B2(n1164), .ZN(n1284)
         );
  XNOR2_X1 U4575 ( .A(n922), .B(n921), .ZN(n914) );
  NAND2_X1 U4576 ( .A1(n921), .A2(n922), .ZN(n918) );
  NAND2_X1 U4577 ( .A1(A2[3]), .A2(n3219), .ZN(n3837) );
  NAND2_X1 U4578 ( .A1(A2[3]), .A2(n3219), .ZN(n3836) );
  OAI221_X1 U4579 ( .B1(reg4[13]), .B2(n2896), .C1(n3676), .C2(n2897), .A(
        n2898), .ZN(n2895) );
  OAI221_X1 U4580 ( .B1(reg4[12]), .B2(n2896), .C1(n3679), .C2(n2897), .A(
        n2898), .ZN(n2799) );
  AOI22_X1 U4581 ( .A1(reg4[11]), .A2(n2897), .B1(n2896), .B2(n3671), .ZN(
        n2924) );
  AOI22_X1 U4582 ( .A1(reg4[10]), .A2(n2897), .B1(n2896), .B2(n3682), .ZN(
        n2946) );
  OAI221_X1 U4583 ( .B1(reg4[8]), .B2(n2896), .C1(n3667), .C2(n2897), .A(n2983), .ZN(n2982) );
  AOI22_X1 U4584 ( .A1(reg4[9]), .A2(n2897), .B1(n2896), .B2(n3681), .ZN(n2966) );
  AOI22_X1 U4585 ( .A1(A2[9]), .A2(n3176), .B1(n3159), .B2(n3158), .ZN(n2854)
         );
  OAI221_X1 U4586 ( .B1(reg4[5]), .B2(n2896), .C1(n3664), .C2(n2897), .A(n3063), .ZN(n3037) );
  OAI221_X1 U4587 ( .B1(reg4[4]), .B2(n2896), .C1(n3668), .C2(n2897), .A(n3083), .ZN(n3060) );
  AOI22_X1 U4588 ( .A1(reg4[0]), .A2(n2897), .B1(n2896), .B2(n3670), .ZN(n3163) );
  AOI22_X1 U4589 ( .A1(reg4[2]), .A2(n2897), .B1(n2896), .B2(n3673), .ZN(n3128) );
  AOI22_X1 U4590 ( .A1(reg4[7]), .A2(n2897), .B1(n2896), .B2(n3672), .ZN(n3012) );
  AOI22_X1 U4591 ( .A1(reg4[1]), .A2(n2897), .B1(n2896), .B2(n3666), .ZN(n3150) );
  AOI22_X1 U4592 ( .A1(reg4[6]), .A2(n2897), .B1(n2896), .B2(n3678), .ZN(n3050) );
  AOI22_X1 U4593 ( .A1(reg4[3]), .A2(n2897), .B1(n2896), .B2(n3665), .ZN(n3109) );
  NAND2_X1 U4594 ( .A1(n2250), .A2(n2251), .ZN(n2247) );
  AOI22_X1 U4595 ( .A1(n1229), .A2(n1230), .B1(n1231), .B2(n1232), .ZN(n1027)
         );
  AOI22_X1 U4596 ( .A1(n1237), .A2(n1238), .B1(n1239), .B2(n1240), .ZN(n1227)
         );
  AOI22_X1 U4597 ( .A1(B0[8]), .A2(n2112), .B1(n2111), .B2(n2005), .ZN(n2242)
         );
  XNOR2_X1 U4598 ( .A(n2691), .B(n2672), .ZN(n2655) );
  OAI221_X1 U4599 ( .B1(B0[6]), .B2(n1874), .C1(n2041), .C2(n1876), .A(n2042), 
        .ZN(n2026) );
  AOI22_X1 U4600 ( .A1(B0[6]), .A2(n1980), .B1(n1979), .B2(n2041), .ZN(n2077)
         );
  AOI22_X1 U4601 ( .A1(B0[6]), .A2(n1988), .B1(n1989), .B2(n2041), .ZN(n2106)
         );
  OAI221_X1 U4602 ( .B1(B0[6]), .B2(n2021), .C1(n2041), .C2(n2022), .A(n2189), 
        .ZN(n2162) );
  AOI22_X1 U4603 ( .A1(B0[6]), .A2(n2006), .B1(n2007), .B2(n2041), .ZN(n2166)
         );
  AOI221_X1 U4604 ( .B1(n1885), .B2(n2041), .C1(n1884), .C2(B0[6]), .A(n2292), 
        .ZN(n2290) );
  AOI22_X1 U4605 ( .A1(B0[6]), .A2(n1997), .B1(n1996), .B2(n2041), .ZN(n2146)
         );
  XNOR2_X1 U4606 ( .A(n2271), .B(n2270), .ZN(n2263) );
  AOI22_X1 U4607 ( .A1(B0[6]), .A2(n2068), .B1(n2067), .B2(n2041), .ZN(n2240)
         );
  AOI22_X1 U4608 ( .A1(B0[6]), .A2(n2148), .B1(n2149), .B2(n2041), .ZN(n2285)
         );
  AOI22_X1 U4609 ( .A1(B2[6]), .A2(n1249), .B1(n1250), .B2(n1142), .ZN(n1385)
         );
  NOR2_X1 U4610 ( .A1(n1504), .A2(n1503), .ZN(p7_C[38]) );
  AOI221_X1 U4611 ( .B1(n529), .B2(B3[9]), .C1(n530), .C2(n654), .A(n655), 
        .ZN(n652) );
  AOI221_X1 U4612 ( .B1(n639), .B2(B3[9]), .C1(n640), .C2(n654), .A(n696), 
        .ZN(n695) );
  AOI22_X1 U4613 ( .A1(B3[9]), .A2(n631), .B1(n630), .B2(n654), .ZN(n670) );
  AOI22_X1 U4614 ( .A1(B3[9]), .A2(n657), .B1(n658), .B2(n654), .ZN(n731) );
  AOI22_X1 U4615 ( .A1(B3[9]), .A2(n648), .B1(n647), .B2(n654), .ZN(n717) );
  OAI221_X1 U4616 ( .B1(B3[9]), .B2(n672), .C1(n654), .C2(n673), .A(n759), 
        .ZN(n736) );
  OAI221_X1 U4617 ( .B1(B3[9]), .B2(n718), .C1(n654), .C2(n719), .A(n819), 
        .ZN(n805) );
  AOI22_X1 U4618 ( .A1(B3[9]), .A2(n732), .B1(n733), .B2(n654), .ZN(n836) );
  OAI221_X1 U4619 ( .B1(B3[9]), .B2(n762), .C1(n654), .C2(n763), .A(n868), 
        .ZN(n867) );
  AOI22_X1 U4620 ( .A1(B3[9]), .A2(n535), .B1(n536), .B2(n654), .ZN(n919) );
  AOI22_X1 U4621 ( .A1(B3[8]), .A2(n527), .B1(n525), .B2(n656), .ZN(n655) );
  AOI22_X1 U4622 ( .A1(B3[8]), .A2(n529), .B1(n530), .B2(n656), .ZN(n669) );
  AOI22_X1 U4623 ( .A1(B3[8]), .A2(n631), .B1(n630), .B2(n656), .ZN(n696) );
  AOI221_X1 U4624 ( .B1(n639), .B2(B3[8]), .C1(n640), .C2(n656), .A(n715), 
        .ZN(n690) );
  OAI221_X1 U4625 ( .B1(B3[8]), .B2(n647), .C1(n656), .C2(n648), .A(n731), 
        .ZN(n730) );
  AOI221_X1 U4626 ( .B1(n657), .B2(B3[8]), .C1(n658), .C2(n656), .A(n765), 
        .ZN(n740) );
  AOI22_X1 U4627 ( .A1(B3[8]), .A2(n673), .B1(n672), .B2(n656), .ZN(n796) );
  OAI221_X1 U4628 ( .B1(B3[8]), .B2(n718), .C1(n656), .C2(n719), .A(n836), 
        .ZN(n826) );
  AOI221_X1 U4629 ( .B1(B3[8]), .B2(n799), .C1(n800), .C2(n656), .A(n889), 
        .ZN(n886) );
  XNOR2_X1 U4630 ( .A(n870), .B(n871), .ZN(n890) );
  AOI22_X1 U4631 ( .A1(B3[8]), .A2(n535), .B1(n536), .B2(n656), .ZN(n935) );
  AOI22_X1 U4632 ( .A1(B3[8]), .A2(n763), .B1(n762), .B2(n656), .ZN(n893) );
  XNOR2_X1 U4633 ( .A(n2870), .B(n2869), .ZN(n2872) );
  XNOR2_X1 U4634 ( .A(n2871), .B(n2872), .ZN(p10_S[34]) );
  AOI22_X1 U4635 ( .A1(B2[3]), .A2(n1123), .B1(n1122), .B2(n3827), .ZN(n1349)
         );
  AOI22_X1 U4636 ( .A1(n2128), .A2(n2129), .B1(n2130), .B2(n2131), .ZN(n1926)
         );
  NAND3_X1 U4637 ( .A1(n2667), .A2(n3839), .A3(n3838), .ZN(n2666) );
  AOI221_X1 U4638 ( .B1(n1428), .B2(B1[5]), .C1(n1429), .C2(n1613), .A(n1624), 
        .ZN(n1603) );
  AOI22_X1 U4639 ( .A1(B1[5]), .A2(n1426), .B1(n1424), .B2(n1613), .ZN(n1612)
         );
  OAI221_X1 U4640 ( .B1(B1[5]), .B2(n1529), .C1(n1613), .C2(n1530), .A(n1656), 
        .ZN(n1642) );
  OAI221_X1 U4641 ( .B1(B1[5]), .B2(n1546), .C1(n1613), .C2(n1547), .A(n1716), 
        .ZN(n1688) );
  AOI22_X1 U4642 ( .A1(B1[5]), .A2(n1556), .B1(n1557), .B2(n1613), .ZN(n1733)
         );
  AOI221_X1 U4643 ( .B1(n1631), .B2(B1[5]), .C1(n1632), .C2(n1613), .A(n1822), 
        .ZN(n1807) );
  XNOR2_X1 U4644 ( .A(n1732), .B(n1741), .ZN(n1763) );
  AOI22_X1 U4645 ( .A1(B2[10]), .A2(n1213), .B1(n1212), .B2(n1092), .ZN(n1289)
         );
  AOI22_X1 U4646 ( .A1(B2[10]), .A2(n1169), .B1(n1168), .B2(n1092), .ZN(n1251)
         );
  AOI22_X1 U4647 ( .A1(B2[10]), .A2(n1182), .B1(n1183), .B2(n1092), .ZN(n1269)
         );
  OAI221_X1 U4648 ( .B1(B2[6]), .B2(n1212), .C1(n1142), .C2(n1213), .A(n1369), 
        .ZN(n1351) );
  XNOR2_X1 U4649 ( .A(n1351), .B(n1350), .ZN(n1356) );
  AOI221_X1 U4650 ( .B1(n1878), .B2(B0[9]), .C1(n1879), .C2(n2003), .A(n2004), 
        .ZN(n2001) );
  AOI221_X1 U4651 ( .B1(n1988), .B2(B0[9]), .C1(n1989), .C2(n2003), .A(n2045), 
        .ZN(n2044) );
  AOI22_X1 U4652 ( .A1(B0[9]), .A2(n2006), .B1(n2007), .B2(n2003), .ZN(n2080)
         );
  OAI221_X1 U4653 ( .B1(B0[9]), .B2(n2021), .C1(n2003), .C2(n2022), .A(n2108), 
        .ZN(n2085) );
  OAI221_X1 U4654 ( .B1(B0[9]), .B2(n2067), .C1(n2003), .C2(n2068), .A(n2168), 
        .ZN(n2154) );
  AOI22_X1 U4655 ( .A1(B0[9]), .A2(n2081), .B1(n2082), .B2(n2003), .ZN(n2185)
         );
  AOI221_X1 U4656 ( .B1(n1878), .B2(B0[5]), .C1(n1879), .C2(n2063), .A(n2074), 
        .ZN(n2053) );
  AOI22_X1 U4657 ( .A1(B0[5]), .A2(n1876), .B1(n1874), .B2(n2063), .ZN(n2062)
         );
  OAI221_X1 U4658 ( .B1(B0[5]), .B2(n1979), .C1(n2063), .C2(n1980), .A(n2106), 
        .ZN(n2092) );
  OAI221_X1 U4659 ( .B1(B0[5]), .B2(n1996), .C1(n2063), .C2(n1997), .A(n2166), 
        .ZN(n2138) );
  AOI22_X1 U4660 ( .A1(B0[5]), .A2(n2006), .B1(n2007), .B2(n2063), .ZN(n2183)
         );
  AOI221_X1 U4661 ( .B1(n2081), .B2(B0[5]), .C1(n2082), .C2(n2063), .A(n2272), 
        .ZN(n2257) );
  AOI22_X1 U4662 ( .A1(B0[5]), .A2(n1884), .B1(n1885), .B2(n2063), .ZN(n2308)
         );
  OAI221_X1 U4663 ( .B1(B0[5]), .B2(n2111), .C1(n2063), .C2(n2112), .A(n2285), 
        .ZN(n2271) );
  AOI22_X1 U4664 ( .A1(B0[5]), .A2(n2068), .B1(n2067), .B2(n2063), .ZN(n2248)
         );
  AOI22_X1 U4665 ( .A1(reg4[3]), .A2(n3047), .B1(n3048), .B2(n3665), .ZN(n3208) );
  AOI22_X1 U4666 ( .A1(A2[13]), .A2(n3841), .B1(n3094), .B2(n2894), .ZN(n3840)
         );
  AOI22_X1 U4667 ( .A1(B1[8]), .A2(n1426), .B1(n1424), .B2(n1555), .ZN(n1554)
         );
  AOI22_X1 U4668 ( .A1(B1[8]), .A2(n1428), .B1(n1429), .B2(n1555), .ZN(n1568)
         );
  AOI22_X1 U4669 ( .A1(B1[8]), .A2(n1530), .B1(n1529), .B2(n1555), .ZN(n1595)
         );
  AOI221_X1 U4670 ( .B1(n1538), .B2(B1[8]), .C1(n1539), .C2(n1555), .A(n1614), 
        .ZN(n1589) );
  OAI221_X1 U4671 ( .B1(B1[8]), .B2(n1546), .C1(n1555), .C2(n1547), .A(n1630), 
        .ZN(n1629) );
  AOI221_X1 U4672 ( .B1(n1556), .B2(B1[8]), .C1(n1557), .C2(n1555), .A(n1664), 
        .ZN(n1639) );
  AOI22_X1 U4673 ( .A1(B1[8]), .A2(n1572), .B1(n1571), .B2(n1555), .ZN(n1695)
         );
  OAI221_X1 U4674 ( .B1(B1[8]), .B2(n1617), .C1(n1555), .C2(n1618), .A(n1735), 
        .ZN(n1725) );
  AOI221_X1 U4675 ( .B1(B1[8]), .B2(n1698), .C1(n1699), .C2(n1555), .A(n1788), 
        .ZN(n1785) );
  XNOR2_X1 U4676 ( .A(n1769), .B(n1770), .ZN(n1789) );
  AOI22_X1 U4677 ( .A1(B1[8]), .A2(n1434), .B1(n1435), .B2(n1555), .ZN(n1834)
         );
  AOI22_X1 U4678 ( .A1(B1[8]), .A2(n1662), .B1(n1661), .B2(n1555), .ZN(n1792)
         );
  AOI22_X1 U4679 ( .A1(B0[10]), .A2(n1876), .B1(n1874), .B2(n1991), .ZN(n1990)
         );
  AOI22_X1 U4680 ( .A1(B0[10]), .A2(n1980), .B1(n1979), .B2(n1991), .ZN(n2008)
         );
  AOI22_X1 U4681 ( .A1(B0[10]), .A2(n1997), .B1(n1996), .B2(n1991), .ZN(n2046)
         );
  AOI22_X1 U4682 ( .A1(B0[10]), .A2(n2022), .B1(n2021), .B2(n1991), .ZN(n2083)
         );
  AOI22_X1 U4683 ( .A1(B0[10]), .A2(n2047), .B1(n2048), .B2(n1991), .ZN(n2108)
         );
  AOI22_X1 U4684 ( .A1(B0[10]), .A2(n2081), .B1(n2082), .B2(n1991), .ZN(n2168)
         );
  AOI22_X1 U4685 ( .A1(B0[10]), .A2(n2068), .B1(n2067), .B2(n1991), .ZN(n2150)
         );
  AOI22_X1 U4686 ( .A1(B0[10]), .A2(n2112), .B1(n2111), .B2(n1991), .ZN(n2188)
         );
  OAI221_X1 U4687 ( .B1(B3[7]), .B2(n525), .C1(n668), .C2(n527), .A(n669), 
        .ZN(n661) );
  AOI22_X1 U4688 ( .A1(B3[7]), .A2(n529), .B1(n530), .B2(n668), .ZN(n693) );
  AOI221_X1 U4689 ( .B1(n639), .B2(B3[7]), .C1(n640), .C2(n668), .A(n728), 
        .ZN(n705) );
  AOI22_X1 U4690 ( .A1(B3[7]), .A2(n631), .B1(n630), .B2(n668), .ZN(n715) );
  AOI22_X1 U4691 ( .A1(B3[7]), .A2(n648), .B1(n647), .B2(n668), .ZN(n765) );
  AOI22_X1 U4692 ( .A1(B3[7]), .A2(n698), .B1(n699), .B2(n668), .ZN(n840) );
  NOR2_X1 U4693 ( .A1(n763), .A2(n668), .ZN(n889) );
  AOI22_X1 U4694 ( .A1(B3[7]), .A2(n673), .B1(n672), .B2(n668), .ZN(n822) );
  AOI22_X1 U4695 ( .A1(B3[7]), .A2(n719), .B1(n718), .B2(n668), .ZN(n865) );
  AOI22_X1 U4696 ( .A1(B3[7]), .A2(n799), .B1(n800), .B2(n668), .ZN(n920) );
  XNOR2_X1 U4697 ( .A(n2219), .B(n2220), .ZN(n2239) );
  AOI222_X1 U4698 ( .A1(n1943), .A2(n1944), .B1(n1943), .B2(n1941), .C1(n1944), 
        .C2(n1941), .ZN(p6_C[41]) );
  XNOR2_X1 U4699 ( .A(n1730), .B(n1766), .ZN(n1732) );
  AOI22_X1 U4700 ( .A1(reg2[10]), .A2(n2601), .B1(n2602), .B2(n3693), .ZN(
        n2667) );
  OAI221_X1 U4701 ( .B1(reg2[13]), .B2(n2471), .C1(n3680), .C2(n3662), .A(
        n2473), .ZN(n2464) );
  OAI221_X1 U4702 ( .B1(reg2[12]), .B2(n2471), .C1(n3690), .C2(n3662), .A(
        n2473), .ZN(n2461) );
  AOI22_X1 U4703 ( .A1(reg2[10]), .A2(n3662), .B1(n2471), .B2(n3693), .ZN(
        n2533) );
  OAI221_X1 U4704 ( .B1(reg2[9]), .B2(n2471), .C1(n3691), .C2(n3662), .A(n2558), .ZN(n2535) );
  AOI22_X1 U4705 ( .A1(reg2[8]), .A2(n3662), .B1(n2471), .B2(n3683), .ZN(n2598) );
  AOI22_X1 U4706 ( .A1(reg2[0]), .A2(n3662), .B1(n2471), .B2(n3689), .ZN(n2752) );
  AOI22_X1 U4707 ( .A1(reg2[2]), .A2(n3662), .B1(n2471), .B2(n3692), .ZN(n2725) );
  AOI22_X1 U4708 ( .A1(reg2[6]), .A2(n3662), .B1(n2471), .B2(n3687), .ZN(n2639) );
  AOI22_X1 U4709 ( .A1(reg2[1]), .A2(n3662), .B1(n2471), .B2(n3684), .ZN(n2734) );
  AOI22_X1 U4710 ( .A1(reg2[7]), .A2(n3662), .B1(n2471), .B2(n3688), .ZN(n2627) );
  OAI221_X1 U4711 ( .B1(reg4[12]), .B2(n2967), .C1(n3679), .C2(n2968), .A(
        n2969), .ZN(n2935) );
  OAI221_X1 U4712 ( .B1(reg4[13]), .B2(n2967), .C1(n3676), .C2(n2968), .A(
        n2969), .ZN(n2950) );
  AOI22_X1 U4713 ( .A1(reg4[11]), .A2(n2968), .B1(n2967), .B2(n3671), .ZN(
        n3011) );
  AOI22_X1 U4714 ( .A1(n3131), .A2(n3132), .B1(n3133), .B2(n3134), .ZN(n3130)
         );
  OAI221_X1 U4715 ( .B1(reg4[0]), .B2(n2967), .C1(n3670), .C2(n2968), .A(n3206), .ZN(n2865) );
  AOI22_X1 U4716 ( .A1(reg4[10]), .A2(n2968), .B1(n2967), .B2(n3682), .ZN(
        n3049) );
  OAI221_X1 U4717 ( .B1(reg4[8]), .B2(n2967), .C1(n3667), .C2(n2968), .A(n3085), .ZN(n3074) );
  AOI22_X1 U4718 ( .A1(reg4[9]), .A2(n2968), .B1(n2967), .B2(n3681), .ZN(n3065) );
  AOI22_X1 U4719 ( .A1(reg4[4]), .A2(n2968), .B1(n2967), .B2(n3668), .ZN(n3170) );
  AOI22_X1 U4720 ( .A1(reg4[3]), .A2(n2968), .B1(n2967), .B2(n3665), .ZN(n3184) );
  AOI22_X1 U4721 ( .A1(reg4[7]), .A2(n2968), .B1(n2967), .B2(n3672), .ZN(n3111) );
  AOI22_X1 U4722 ( .A1(reg4[2]), .A2(n2968), .B1(n2967), .B2(n3673), .ZN(n3195) );
  AOI22_X1 U4723 ( .A1(reg4[6]), .A2(n2968), .B1(n2967), .B2(n3678), .ZN(n3138) );
  AOI22_X1 U4724 ( .A1(reg4[1]), .A2(n2968), .B1(n2967), .B2(n3666), .ZN(n3201) );
  AOI22_X1 U4725 ( .A1(reg4[5]), .A2(n2968), .B1(n2967), .B2(n3664), .ZN(n3146) );
  AOI22_X1 U4726 ( .A1(B2[9]), .A2(n985), .B1(n986), .B2(n1104), .ZN(n1368) );
  AOI22_X1 U4727 ( .A1(B2[9]), .A2(n1182), .B1(n1183), .B2(n1104), .ZN(n1286)
         );
  OAI221_X1 U4728 ( .B1(B2[9]), .B2(n1168), .C1(n1104), .C2(n1169), .A(n1269), 
        .ZN(n1255) );
  OAI221_X1 U4729 ( .B1(B0[2]), .B2(n1874), .C1(n2133), .C2(n1876), .A(n2134), 
        .ZN(n2121) );
  AOI22_X1 U4730 ( .A1(B0[2]), .A2(n1980), .B1(n1979), .B2(n2133), .ZN(n2190)
         );
  AOI22_X1 U4731 ( .A1(B0[2]), .A2(n1997), .B1(n1996), .B2(n2133), .ZN(n2230)
         );
  AOI22_X1 U4732 ( .A1(B0[2]), .A2(n2022), .B1(n2021), .B2(n2133), .ZN(n2273)
         );
  AOI22_X1 U4733 ( .A1(B0[2]), .A2(n2068), .B1(n2067), .B2(n2133), .ZN(n2295)
         );
  AOI22_X1 U4734 ( .A1(B0[2]), .A2(n2081), .B1(n2082), .B2(n2133), .ZN(n2302)
         );
  AOI22_X1 U4735 ( .A1(B0[2]), .A2(n2148), .B1(n2149), .B2(n2133), .ZN(n2311)
         );
  NOR2_X1 U4736 ( .A1(n2404), .A2(n2403), .ZN(p11_C[38]) );
  AOI22_X1 U4737 ( .A1(B2[7]), .A2(n1249), .B1(n1250), .B2(n1118), .ZN(n1369)
         );
  AOI22_X1 U4738 ( .A1(B2[7]), .A2(n1169), .B1(n1168), .B2(n1118), .ZN(n1313)
         );
  AOI22_X1 U4739 ( .A1(B2[7]), .A2(n1123), .B1(n1122), .B2(n1118), .ZN(n1272)
         );
  NOR2_X1 U4740 ( .A1(n1213), .A2(n1118), .ZN(n1338) );
  AOI22_X1 U4741 ( .A1(A1[9]), .A2(n2730), .B1(n2713), .B2(n2712), .ZN(n2404)
         );
  AOI22_X1 U4742 ( .A1(B1[10]), .A2(n1662), .B1(n1661), .B2(n1541), .ZN(n1738)
         );
  AOI221_X1 U4743 ( .B1(n1435), .B2(n1541), .C1(n1434), .C2(B1[10]), .A(n1787), 
        .ZN(n1786) );
  AOI22_X1 U4744 ( .A1(B1[10]), .A2(n1618), .B1(n1617), .B2(n1541), .ZN(n1700)
         );
  AOI22_X1 U4745 ( .A1(B1[10]), .A2(n1631), .B1(n1632), .B2(n1541), .ZN(n1718)
         );
  OAI221_X1 U4746 ( .B1(B0[7]), .B2(n1874), .C1(n2017), .C2(n1876), .A(n2018), 
        .ZN(n2010) );
  AOI22_X1 U4747 ( .A1(B0[7]), .A2(n1878), .B1(n1879), .B2(n2017), .ZN(n2042)
         );
  AOI221_X1 U4748 ( .B1(n1988), .B2(B0[7]), .C1(n1989), .C2(n2017), .A(n2077), 
        .ZN(n2054) );
  AOI22_X1 U4749 ( .A1(B0[7]), .A2(n1980), .B1(n1979), .B2(n2017), .ZN(n2064)
         );
  AOI22_X1 U4750 ( .A1(B0[7]), .A2(n1997), .B1(n1996), .B2(n2017), .ZN(n2114)
         );
  AOI22_X1 U4751 ( .A1(B0[7]), .A2(n2047), .B1(n2048), .B2(n2017), .ZN(n2189)
         );
  NOR2_X1 U4752 ( .A1(n2112), .A2(n2017), .ZN(n2238) );
  AOI22_X1 U4753 ( .A1(B0[7]), .A2(n2022), .B1(n2021), .B2(n2017), .ZN(n2171)
         );
  AOI22_X1 U4754 ( .A1(B0[7]), .A2(n2068), .B1(n2067), .B2(n2017), .ZN(n2214)
         );
  XNOR2_X1 U4755 ( .A(n1505), .B(n1506), .ZN(p7_S[37]) );
  AOI221_X1 U4756 ( .B1(n1698), .B2(B1[3]), .C1(n1699), .C2(n1665), .A(n1859), 
        .ZN(n1849) );
  OAI22_X1 U4757 ( .A1(n1849), .A2(n1850), .B1(n1851), .B2(n3714), .ZN(
        p7_C[36]) );
  AOI222_X1 U4758 ( .A1(n1501), .A2(n1502), .B1(n1501), .B2(n1499), .C1(n1502), 
        .C2(n1499), .ZN(p7_C[39]) );
  AOI22_X1 U4759 ( .A1(B1[5]), .A2(n1572), .B1(n1571), .B2(n1613), .ZN(n1765)
         );
  AOI22_X1 U4760 ( .A1(B1[5]), .A2(n1618), .B1(n1617), .B2(n1613), .ZN(n1798)
         );
  AOI22_X1 U4761 ( .A1(B1[5]), .A2(n1434), .B1(n1435), .B2(n1613), .ZN(n1858)
         );
  OAI221_X1 U4762 ( .B1(B1[5]), .B2(n1661), .C1(n1613), .C2(n1662), .A(n1835), 
        .ZN(n1821) );
  XNOR2_X1 U4763 ( .A(n2634), .B(n2666), .ZN(n2636) );
  XNOR2_X1 U4764 ( .A(n1056), .B(n1057), .ZN(p8_S[37]) );
  XNOR2_X1 U4765 ( .A(n2399), .B(n2400), .ZN(p11_S[39]) );
  AOI22_X1 U4766 ( .A1(reg2[7]), .A2(n2601), .B1(n2602), .B2(n3688), .ZN(n2721) );
  OAI221_X1 U4767 ( .B1(B1[9]), .B2(n1661), .C1(n1553), .C2(n1662), .A(n1767), 
        .ZN(n1766) );
  AOI22_X1 U4768 ( .A1(B1[10]), .A2(n1698), .B1(n1699), .B2(n1541), .ZN(n1767)
         );
  XNOR2_X1 U4769 ( .A(n1517), .B(n1518), .ZN(n1516) );
  OAI211_X1 U4770 ( .C1(n1517), .C2(n1515), .A(n1520), .B(n1519), .ZN(n1855)
         );
  NAND2_X1 U4771 ( .A1(n1517), .A2(n1515), .ZN(n1856) );
  AOI221_X1 U4772 ( .B1(n529), .B2(B3[5]), .C1(n530), .C2(n714), .A(n725), 
        .ZN(n704) );
  AOI22_X1 U4773 ( .A1(B3[5]), .A2(n527), .B1(n525), .B2(n714), .ZN(n713) );
  OAI221_X1 U4774 ( .B1(B3[5]), .B2(n630), .C1(n714), .C2(n631), .A(n757), 
        .ZN(n743) );
  OAI221_X1 U4775 ( .B1(B3[5]), .B2(n647), .C1(n714), .C2(n648), .A(n817), 
        .ZN(n789) );
  AOI22_X1 U4776 ( .A1(B3[5]), .A2(n657), .B1(n658), .B2(n714), .ZN(n834) );
  AOI221_X1 U4777 ( .B1(n698), .B2(B3[5]), .C1(n699), .C2(n714), .A(n882), 
        .ZN(n854) );
  AOI221_X1 U4778 ( .B1(n732), .B2(B3[5]), .C1(n733), .C2(n714), .A(n923), 
        .ZN(n908) );
  OAI221_X1 U4779 ( .B1(B3[5]), .B2(n762), .C1(n714), .C2(n763), .A(n936), 
        .ZN(n922) );
  AOI22_X1 U4780 ( .A1(B3[5]), .A2(n535), .B1(n536), .B2(n714), .ZN(n959) );
  AOI22_X1 U4781 ( .A1(B3[5]), .A2(n719), .B1(n718), .B2(n714), .ZN(n899) );
  AOI22_X1 U4782 ( .A1(B3[5]), .A2(n673), .B1(n672), .B2(n714), .ZN(n866) );
  AOI22_X1 U4783 ( .A1(B3[10]), .A2(n527), .B1(n525), .B2(n642), .ZN(n641) );
  AOI22_X1 U4784 ( .A1(B3[10]), .A2(n631), .B1(n630), .B2(n642), .ZN(n659) );
  AOI221_X1 U4785 ( .B1(n639), .B2(B3[10]), .C1(n640), .C2(n642), .A(n670), 
        .ZN(n664) );
  AOI22_X1 U4786 ( .A1(B3[10]), .A2(n648), .B1(n647), .B2(n642), .ZN(n697) );
  AOI221_X1 U4787 ( .B1(n657), .B2(B3[10]), .C1(n658), .C2(n642), .A(n717), 
        .ZN(n703) );
  AOI22_X1 U4788 ( .A1(B3[10]), .A2(n673), .B1(n672), .B2(n642), .ZN(n734) );
  AOI22_X1 U4789 ( .A1(B3[10]), .A2(n698), .B1(n699), .B2(n642), .ZN(n759) );
  AOI22_X1 U4790 ( .A1(B3[10]), .A2(n732), .B1(n733), .B2(n642), .ZN(n819) );
  AOI22_X1 U4791 ( .A1(B3[10]), .A2(n719), .B1(n718), .B2(n642), .ZN(n801) );
  AOI22_X1 U4792 ( .A1(B3[10]), .A2(n763), .B1(n762), .B2(n642), .ZN(n839) );
  XNOR2_X1 U4793 ( .A(n831), .B(n867), .ZN(n833) );
  AOI22_X1 U4794 ( .A1(B3[10]), .A2(n799), .B1(n800), .B2(n642), .ZN(n868) );
  XNOR2_X1 U4795 ( .A(n606), .B(n607), .ZN(p9_S[37]) );
  XNOR2_X1 U4796 ( .A(n2421), .B(n2422), .ZN(p11_S[34]) );
  NOR3_X1 U4797 ( .A1(n3842), .A2(n3843), .A3(n3115), .ZN(n3090) );
  AOI222_X1 U4798 ( .A1(n2794), .A2(n2882), .B1(n2794), .B2(n2796), .C1(n2882), 
        .C2(n2796), .ZN(p10_C[53]) );
  XNOR2_X1 U4799 ( .A(n2790), .B(n2791), .ZN(p10_S[54]) );
  XNOR2_X1 U4800 ( .A(n3149), .B(n3148), .ZN(n3154) );
  AOI222_X1 U4801 ( .A1(n2851), .A2(n2852), .B1(n2851), .B2(n2849), .C1(n2852), 
        .C2(n2849), .ZN(p10_C[39]) );
  AOI22_X1 U4802 ( .A1(B2[5]), .A2(n1169), .B1(n1168), .B2(n1164), .ZN(n1348)
         );
  AOI22_X1 U4803 ( .A1(B2[5]), .A2(n985), .B1(n986), .B2(n1164), .ZN(n1408) );
  OAI221_X1 U4804 ( .B1(B2[5]), .B2(n1212), .C1(n1164), .C2(n1213), .A(n1385), 
        .ZN(n1371) );
  AOI222_X1 U4805 ( .A1(n2397), .A2(n2398), .B1(n2397), .B2(n2395), .C1(n2398), 
        .C2(n2395), .ZN(p11_C[40]) );
  XNOR2_X1 U4806 ( .A(n2395), .B(n2396), .ZN(p11_S[40]) );
  XNOR2_X1 U4807 ( .A(n618), .B(n619), .ZN(n617) );
  XNOR2_X1 U4808 ( .A(n2703), .B(n2702), .ZN(n2708) );
  XNOR2_X1 U4809 ( .A(n3105), .B(n3095), .ZN(n3094) );
  XNOR2_X1 U4810 ( .A(n3124), .B(n3125), .ZN(n3142) );
  NAND2_X1 U4811 ( .A1(n2648), .A2(n2444), .ZN(n3845) );
  XNOR2_X1 U4812 ( .A(n1955), .B(n1956), .ZN(p6_S[37]) );
  AOI222_X1 U4813 ( .A1(n1892), .A2(n1893), .B1(n1892), .B2(n1891), .C1(n1893), 
        .C2(n1891), .ZN(p6_C[54]) );
  XNOR2_X1 U4814 ( .A(n2636), .B(n2644), .ZN(n2664) );
  NAND2_X1 U4815 ( .A1(n2753), .A2(n2754), .ZN(p11_C[36]) );
  AOI22_X1 U4816 ( .A1(B2[2]), .A2(n1081), .B1(n1080), .B2(n1234), .ZN(n1291)
         );
  NAND2_X1 U4817 ( .A1(n1068), .A2(n1066), .ZN(n1406) );
  OAI211_X1 U4818 ( .C1(n1068), .C2(n1066), .A(n1071), .B(n1070), .ZN(n1405)
         );
  AOI22_X1 U4819 ( .A1(B2[2]), .A2(n1098), .B1(n1097), .B2(n1234), .ZN(n1330)
         );
  XNOR2_X1 U4820 ( .A(n1068), .B(n1069), .ZN(n1067) );
  AOI22_X1 U4821 ( .A1(B2[2]), .A2(n1123), .B1(n1122), .B2(n1234), .ZN(n1373)
         );
  AOI22_X1 U4822 ( .A1(B2[2]), .A2(n1169), .B1(n1168), .B2(n1234), .ZN(n1395)
         );
  AOI22_X1 U4823 ( .A1(B2[2]), .A2(n1182), .B1(n1183), .B2(n1234), .ZN(n1402)
         );
  AOI22_X1 U4824 ( .A1(B2[2]), .A2(n1249), .B1(n1250), .B2(n1234), .ZN(n1411)
         );
  AOI22_X1 U4825 ( .A1(B2[2]), .A2(n985), .B1(n986), .B2(n1234), .ZN(n1418) );
  AOI22_X1 U4826 ( .A1(B2[2]), .A2(n1213), .B1(n1212), .B2(n1234), .ZN(n1409)
         );
  NAND2_X1 U4827 ( .A1(n1967), .A2(n1965), .ZN(n2306) );
  OAI211_X1 U4828 ( .C1(n1967), .C2(n1965), .A(n1970), .B(n1969), .ZN(n2305)
         );
  AOI222_X1 U4829 ( .A1(n2874), .A2(n2873), .B1(n2874), .B2(n2872), .C1(n2873), 
        .C2(n2872), .ZN(p10_C[34]) );
  NOR2_X1 U4830 ( .A1(n2854), .A2(n2853), .ZN(p10_C[38]) );
  OAI221_X1 U4831 ( .B1(reg2[13]), .B2(n2561), .C1(n3680), .C2(n2562), .A(
        n2563), .ZN(n2537) );
  OAI221_X1 U4832 ( .B1(reg2[12]), .B2(n2561), .C1(n3690), .C2(n2562), .A(
        n2563), .ZN(n2545) );
  NOR2_X1 U4833 ( .A1(n2428), .A2(n2427), .ZN(p11_C[32]) );
  OAI221_X1 U4834 ( .B1(reg2[11]), .B2(n2561), .C1(n3686), .C2(n2562), .A(
        n2624), .ZN(n2623) );
  AOI22_X1 U4835 ( .A1(reg2[10]), .A2(n2562), .B1(n2561), .B2(n3693), .ZN(
        n2643) );
  OAI221_X1 U4836 ( .B1(reg2[5]), .B2(n2561), .C1(n3677), .C2(n2562), .A(n2737), .ZN(n2723) );
  AOI22_X1 U4837 ( .A1(reg2[8]), .A2(n2562), .B1(n2561), .B2(n3683), .ZN(n2694) );
  AOI22_X1 U4838 ( .A1(reg2[4]), .A2(n2562), .B1(n2561), .B2(n3685), .ZN(n2751) );
  OAI221_X1 U4839 ( .B1(reg2[2]), .B2(n2561), .C1(n3692), .C2(n2562), .A(n2762), .ZN(n2414) );
  AOI22_X1 U4840 ( .A1(reg2[0]), .A2(n2562), .B1(n2561), .B2(n3689), .ZN(n2769) );
  OAI221_X1 U4841 ( .B1(reg2[1]), .B2(n2561), .C1(n3684), .C2(n2562), .A(n2763), .ZN(n2419) );
  XNOR2_X1 U4842 ( .A(n2849), .B(n2850), .ZN(p10_S[39]) );
  OAI221_X1 U4843 ( .B1(B3[2]), .B2(n525), .C1(n784), .C2(n527), .A(n785), 
        .ZN(n772) );
  AOI22_X1 U4844 ( .A1(B3[2]), .A2(n631), .B1(n630), .B2(n784), .ZN(n841) );
  AOI22_X1 U4845 ( .A1(B3[2]), .A2(n648), .B1(n647), .B2(n784), .ZN(n881) );
  AOI22_X1 U4846 ( .A1(B3[2]), .A2(n673), .B1(n672), .B2(n784), .ZN(n924) );
  AOI22_X1 U4847 ( .A1(B3[2]), .A2(n719), .B1(n718), .B2(n784), .ZN(n946) );
  AOI22_X1 U4848 ( .A1(B3[2]), .A2(n732), .B1(n733), .B2(n784), .ZN(n953) );
  AOI22_X1 U4849 ( .A1(B3[2]), .A2(n799), .B1(n800), .B2(n784), .ZN(n962) );
  AOI22_X1 U4850 ( .A1(B3[2]), .A2(n763), .B1(n762), .B2(n784), .ZN(n960) );
  AOI22_X1 U4851 ( .A1(B3[2]), .A2(n535), .B1(n536), .B2(n784), .ZN(n969) );
  OAI221_X1 U4852 ( .B1(B1[2]), .B2(n1424), .C1(n1683), .C2(n1426), .A(n1684), 
        .ZN(n1671) );
  AOI22_X1 U4853 ( .A1(B1[2]), .A2(n1530), .B1(n1529), .B2(n1683), .ZN(n1740)
         );
  AOI22_X1 U4854 ( .A1(B1[2]), .A2(n1547), .B1(n1546), .B2(n1683), .ZN(n1780)
         );
  AOI22_X1 U4855 ( .A1(B1[2]), .A2(n1572), .B1(n1571), .B2(n1683), .ZN(n1823)
         );
  AOI22_X1 U4856 ( .A1(B1[2]), .A2(n1618), .B1(n1617), .B2(n1683), .ZN(n1845)
         );
  AOI22_X1 U4857 ( .A1(B1[2]), .A2(n1631), .B1(n1632), .B2(n1683), .ZN(n1852)
         );
  AOI22_X1 U4858 ( .A1(B1[2]), .A2(n1698), .B1(n1699), .B2(n1683), .ZN(n1861)
         );
  AOI22_X1 U4859 ( .A1(B1[2]), .A2(n1662), .B1(n1661), .B2(n1683), .ZN(n1859)
         );
  AOI22_X1 U4860 ( .A1(B1[2]), .A2(n1434), .B1(n1435), .B2(n1683), .ZN(n1868)
         );
  OAI221_X1 U4861 ( .B1(reg4[13]), .B2(n2921), .C1(n3676), .C2(n2922), .A(
        n2923), .ZN(n2914) );
  OAI221_X1 U4862 ( .B1(reg4[12]), .B2(n2921), .C1(n3679), .C2(n2922), .A(
        n2923), .ZN(n2911) );
  AOI22_X1 U4863 ( .A1(reg4[10]), .A2(n2922), .B1(n2921), .B2(n3682), .ZN(
        n2986) );
  AOI22_X1 U4864 ( .A1(reg4[11]), .A2(n2922), .B1(n2921), .B2(n3671), .ZN(
        n2970) );
  OAI221_X1 U4865 ( .B1(reg4[6]), .B2(n2921), .C1(n3678), .C2(n2922), .A(n3089), .ZN(n3059) );
  AOI22_X1 U4866 ( .A1(reg4[7]), .A2(n2922), .B1(n2921), .B2(n3672), .ZN(n3070) );
  AOI22_X1 U4867 ( .A1(reg4[2]), .A2(n2922), .B1(n2921), .B2(n3673), .ZN(n3171) );
  XNOR2_X1 U4868 ( .A(n3090), .B(n3082), .ZN(n3110) );
  AOI22_X1 U4869 ( .A1(reg4[1]), .A2(n2922), .B1(n2921), .B2(n3666), .ZN(n3180) );
  AOI22_X1 U4870 ( .A1(reg4[3]), .A2(n2922), .B1(n2921), .B2(n3665), .ZN(n3147) );
  AOI22_X1 U4871 ( .A1(reg4[5]), .A2(n2922), .B1(n2921), .B2(n3664), .ZN(n3115) );
  OAI221_X1 U4872 ( .B1(reg2[12]), .B2(n2517), .C1(n3690), .C2(n3826), .A(
        n2519), .ZN(n2485) );
  OAI221_X1 U4873 ( .B1(reg2[13]), .B2(n2517), .C1(n3680), .C2(n3826), .A(
        n2519), .ZN(n2500) );
  OAI221_X1 U4874 ( .B1(reg2[11]), .B2(n2517), .C1(n3686), .C2(n3826), .A(
        n2560), .ZN(n2559) );
  AOI22_X1 U4875 ( .A1(reg2[10]), .A2(n3826), .B1(n2517), .B2(n3693), .ZN(
        n2603) );
  AOI22_X1 U4876 ( .A1(reg2[9]), .A2(n3826), .B1(n2517), .B2(n3691), .ZN(n2622) );
  OAI221_X1 U4877 ( .B1(reg2[0]), .B2(n2517), .C1(n3689), .C2(n3826), .A(n2760), .ZN(n2415) );
  AOI22_X1 U4878 ( .A1(reg2[8]), .A2(n3826), .B1(n2517), .B2(n3683), .ZN(n2640) );
  AOI22_X1 U4879 ( .A1(reg2[4]), .A2(n3826), .B1(n2517), .B2(n3685), .ZN(n2724) );
  AOI22_X1 U4880 ( .A1(reg2[6]), .A2(n3826), .B1(n2517), .B2(n3687), .ZN(n2692) );
  AOI22_X1 U4881 ( .A1(reg2[3]), .A2(n3826), .B1(n2517), .B2(n3669), .ZN(n2738) );
  AOI22_X1 U4882 ( .A1(reg2[2]), .A2(n3826), .B1(n2517), .B2(n3692), .ZN(n2749) );
  AOI22_X1 U4883 ( .A1(reg2[5]), .A2(n3826), .B1(n2517), .B2(n3677), .ZN(n2700) );
  AOI22_X1 U4884 ( .A1(reg2[1]), .A2(n3826), .B1(n2517), .B2(n3684), .ZN(n2755) );
  OAI221_X1 U4885 ( .B1(reg4[13]), .B2(n3836), .C1(n3676), .C2(n3009), .A(
        n3010), .ZN(n2980) );
  OAI221_X1 U4886 ( .B1(reg4[12]), .B2(n3837), .C1(n3679), .C2(n3009), .A(
        n3010), .ZN(n2994) );
  OAI221_X1 U4887 ( .B1(reg4[11]), .B2(n3837), .C1(n3671), .C2(n3009), .A(
        n3067), .ZN(n3066) );
  OAI22_X1 U4888 ( .A1(reg4[9]), .A2(n2782), .B1(reg4[7]), .B2(n3836), .ZN(
        n3135) );
  AOI22_X1 U4889 ( .A1(reg4[10]), .A2(n3009), .B1(n3836), .B2(n3682), .ZN(
        n3088) );
  NOR2_X1 U4890 ( .A1(n2878), .A2(n2877), .ZN(p10_C[32]) );
  OAI221_X1 U4891 ( .B1(reg4[5]), .B2(n3837), .C1(n3664), .C2(n3009), .A(n3183), .ZN(n3169) );
  AOI22_X1 U4892 ( .A1(reg4[8]), .A2(n3009), .B1(n3836), .B2(n3667), .ZN(n3140) );
  OAI221_X1 U4893 ( .B1(reg4[6]), .B2(n3836), .C1(n3678), .C2(n3009), .A(n3167), .ZN(n3149) );
  AOI22_X1 U4894 ( .A1(reg4[4]), .A2(n3009), .B1(n3837), .B2(n3668), .ZN(n3197) );
  OAI221_X1 U4895 ( .B1(reg4[2]), .B2(n3837), .C1(n3673), .C2(n3009), .A(n3208), .ZN(n2864) );
  AOI22_X1 U4896 ( .A1(reg4[0]), .A2(n3009), .B1(n3836), .B2(n3670), .ZN(n3216) );
  OAI221_X1 U4897 ( .B1(reg4[1]), .B2(n3837), .C1(n3666), .C2(n3009), .A(n3209), .ZN(n2869) );
endmodule

